netcdf bigdata {
// Test file containing decent amount of real data. Not huge, but hopefully
// enough to provide a meaningful test of data variable creation.

dimensions:
	height = 1 ;
	latitude = 73 ;
	longitude = 96 ;
	time = 1 ;

variables:
	float height(height) ;
		height:units = "m" ;
		height:axis = "Z" ;
		height:standard_name = "height" ;
	float latitude(latitude) ;
		latitude:units = "degrees_north" ;
		latitude:axis = "Y" ;
		latitude:standard_name = "latitude" ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
	float tas(time, height, latitude, longitude) ;
		tas:_FillValue = -1.0e30f ;
		tas:long_name = "Temperature at 1.5 m" ;
		tas:units = "K" ;
		tas:standard_name = "air_temperature" ;
		tas:cell_methods = "time: mean" ;
	float time(time) ;
		time:units = "days since 1960-1-1" ;
		time:calendar = "360_day" ;
		time:axis = "T" ;
		time:standard_name = "time" ;

// global attributes:
		:Conventions = "CF-1.0" ;

data:

 time = 5730 ;

 height = 1.5 ;

 latitude = 90, 87.5, 85, 82.5, 80, 77.5, 75, 72.5, 70, 67.5, 65, 62.5, 60, 
    57.5, 55, 52.5, 50, 47.5, 45, 42.5, 40, 37.5, 35, 32.5, 30, 27.5, 25, 
    22.5, 20, 17.5, 15, 12.5, 10, 7.5, 5, 2.5, 0, -2.5, -5, -7.5, -10, -12.5, 
    -15, -17.5, -20, -22.5, -25, -27.5, -30, -32.5, -35, -37.5, -40, -42.5, 
    -45, -47.5, -50, -52.5, -55, -57.5, -60, -62.5, -65, -67.5, -70, -72.5, 
    -75, -77.5, -80, -82.5, -85, -87.5, -90 ;

 longitude = 0, 3.75, 7.5, 11.25, 15, 18.75, 22.5, 26.25, 30, 33.75, 37.5, 
    41.25, 45, 48.75, 52.5, 56.25, 60, 63.75, 67.5, 71.25, 75, 78.75, 82.5, 
    86.25, 90, 93.75, 97.5, 101.25, 105, 108.75, 112.5, 116.25, 120, 123.75, 
    127.5, 131.25, 135, 138.75, 142.5, 146.25, 150, 153.75, 157.5, 161.25, 
    165, 168.75, 172.5, 176.25, 180, 183.75, 187.5, 191.25, 195, 198.75, 
    202.5, 206.25, 210, 213.75, 217.5, 221.25, 225, 228.75, 232.5, 236.25, 
    240, 243.75, 247.5, 251.25, 255, 258.75, 262.5, 266.25, 270, 273.75, 
    277.5, 281.25, 285, 288.75, 292.5, 296.25, 300, 303.75, 307.5, 311.25, 
    315, 318.75, 322.5, 326.25, 330, 333.75, 337.5, 341.25, 345, 348.75, 
    352.5, 356.25 ;

 tas =
  253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 
    253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 
    253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 
    253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 
    253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 
    253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 
    253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 
    253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 
    253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 
    253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 
    253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 
    253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 
    253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 253.9404, 
    253.9404, 253.9404, 253.9404, 253.9404, 253.9404,
  254.3543, 254.2611, 254.1507, 254.1776, 254.254, 254.3674, 254.4031, 
    254.3733, 254.369, 254.3443, 254.2977, 254.2474, 254.2255, 254.2256, 
    254.2469, 254.2354, 254.2704, 254.3251, 254.2975, 254.3239, 254.3504, 
    254.3737, 254.4019, 254.398, 254.3861, 254.4079, 254.4458, 254.4165, 
    254.4385, 254.5314, 254.4496, 254.4688, 254.4838, 254.4405, 254.3126, 
    254.1913, 254.1905, 254.3424, 254.1043, 253.9902, 253.9785, 253.9292, 
    253.926, 253.94, 253.9092, 253.903, 253.9057, 253.924, 253.9212, 
    253.8814, 253.8538, 253.8013, 253.7387, 253.6775, 253.5729, 253.4217, 
    253.3818, 253.2512, 253.1728, 253.1, 253.0269, 252.9453, 252.9362, 
    252.9555, 252.9277, 252.8815, 252.9186, 252.9474, 252.9958, 253.0928, 
    253.1926, 253.3568, 253.4521, 253.7956, 254.2065, 253.641, 253.4, 
    253.4077, 253.7732, 254.1251, 253.6547, 253.4639, 253.6717, 253.7958, 
    253.776, 253.9323, 254.141, 254.3075, 254.3876, 254.526, 254.5332, 
    254.2091, 254.1118, 254.1713, 254.2375, 254.3057,
  257.4072, 257.6165, 257.6294, 257.4802, 257.3813, 257.3755, 257.2991, 
    257.1636, 257.1077, 257.0017, 256.9089, 256.7175, 256.5659, 256.4578, 
    256.365, 256.1895, 256.0889, 256.1313, 256.0698, 256.1216, 256.135, 
    256.1846, 256.1973, 256.2202, 256.2803, 256.2886, 256.3484, 256.2083, 
    256.1519, 256.1799, 256.1174, 256.0981, 255.9859, 255.7801, 255.5427, 
    255.3197, 255.1875, 255.0418, 254.8577, 254.6478, 254.4525, 254.3221, 
    254.192, 254.0809, 253.9526, 253.8475, 253.7396, 253.6752, 253.5763, 
    253.4936, 253.4174, 253.3372, 253.2603, 253.1582, 253.0581, 252.9474, 
    252.899, 252.8426, 252.829, 252.8388, 252.9102, 252.9695, 253.1409, 
    253.2245, 253.2737, 253.159, 253.0922, 252.9199, 252.8014, 252.6801, 
    252.9003, 253.29, 253.4745, 254.1756, 255.2845, 253.2831, 252.7031, 
    252.7956, 253.8406, 255.5837, 254.3174, 254.2974, 254.6771, 254.2766, 
    253.2596, 253.7035, 254.0449, 254.4254, 254.6255, 255.5531, 256.6099, 
    255.8641, 255.8233, 256.0066, 256.364, 256.918,
  262.0264, 263.2991, 263.811, 263.2476, 262.5359, 261.9282, 261.4797, 
    261.114, 260.856, 260.5352, 260.1841, 259.8684, 259.4243, 259.1433, 
    258.8525, 258.282, 257.8135, 257.7964, 257.4829, 257.4849, 257.5718, 
    257.6497, 257.5618, 257.5996, 258.1897, 258.1179, 258.3892, 257.718, 
    257.6335, 257.6497, 257.4766, 257.4873, 257.3208, 257.0635, 256.7629, 
    256.4363, 256.2041, 255.956, 255.642, 255.3229, 255.0573, 254.878, 
    254.6859, 254.4581, 254.2936, 254.1652, 254.0236, 253.9018, 253.8038, 
    253.7044, 253.5996, 253.4953, 253.3872, 253.273, 253.1831, 253.1211, 
    253.0689, 253.0358, 253.0595, 253.1864, 253.3685, 253.6092, 253.8512, 
    253.9689, 254.022, 253.9802, 253.8749, 253.6406, 253.3695, 253.3193, 
    254.0359, 255.4691, 254.2907, 254.8341, 257.1116, 245.2807, 245.762, 
    246.8125, 250.6811, 257.1191, 255.9059, 255.6642, 256.4453, 257.2129, 
    248.985, 248.9404, 248.8404, 249.8711, 253.2409, 254.5551, 256.8752, 
    256.0781, 256.4971, 257.2009, 258.1777, 260.0786,
  267.6328, 269.623, 271.1628, 271.4504, 270.7388, 269.8381, 269.4402, 
    268.8076, 267.7957, 266.4897, 265.6897, 265.0435, 264.1416, 263.0354, 
    261.804, 260.6838, 259.916, 259.6748, 259.3147, 259.3765, 259.6948, 
    259.3027, 258.6753, 258.7092, 258.9153, 258.9407, 258.645, 258.0063, 
    258.2134, 259.1316, 258.9036, 258.8381, 258.2932, 257.9016, 257.6045, 
    257.218, 257.0071, 256.7947, 256.4636, 256.1118, 255.8492, 255.6378, 
    255.3848, 255.0385, 254.8974, 254.8079, 254.6638, 254.4797, 254.2798, 
    254.0724, 253.8681, 253.666, 253.5434, 253.5275, 253.5311, 253.5612, 
    253.5034, 253.4038, 253.3349, 253.3392, 253.4588, 253.7309, 254.1948, 
    254.6292, 255.103, 255.4667, 255.6585, 255.5991, 255.3445, 255.3411, 
    256.064, 258.2991, 248.1934, 251.0074, 250.2355, 247.1958, 247.1451, 
    248.5587, 252.3189, 252.6819, 249.2516, 249.3124, 248.8176, 248.1108, 
    247.2557, 247.0659, 247.7768, 249.6517, 251.6351, 252.5743, 253.3398, 
    254.1905, 258.2263, 259.1633, 261.2957, 264.6111,
  269.7473, 271.469, 272.9893, 273.7878, 272.6621, 271.1653, 270.9409, 
    271.1394, 270.644, 269.0776, 267.5764, 266.501, 265.4436, 264.2773, 
    263.0974, 262.2812, 261.5847, 261.1216, 260.7041, 260.4734, 260.7988, 
    260.1609, 259.4858, 259.5591, 259.1638, 259.4475, 259.8992, 254.4664, 
    254.7238, 259.8833, 260.1123, 260.4075, 259.1799, 258.7563, 258.8486, 
    258.7583, 258.5325, 258.4329, 258.3765, 258.1719, 257.938, 257.6165, 
    257.0659, 256.3689, 256.042, 255.8509, 255.6032, 255.3233, 255.1177, 
    254.9402, 254.7587, 254.4346, 254.1779, 254.1844, 254.0645, 254.1862, 
    254.2216, 254.1133, 253.9974, 253.9, 253.8423, 254.0931, 254.7911, 
    255.2418, 255.872, 256.3738, 256.5388, 256.6538, 256.5913, 256.8896, 
    257.6934, 258.7744, 251.4213, 251.5077, 250.1868, 249.0246, 261.5503, 
    263.5845, 248.8973, 251.1168, 251.2307, 250.9926, 249.1111, 246.5075, 
    244.6142, 243.9779, 244.4057, 246.4378, 249.5846, 251.9405, 253.3135, 
    260.521, 260.2122, 261.6831, 264.4133, 267.4282,
  272.2593, 273.2273, 274.2837, 275.3621, 275.8113, 274.5054, 273.3176, 
    273.3711, 272.4373, 270.0396, 268.0854, 266.4429, 265.1311, 264.1973, 
    263.2505, 262.3931, 261.7888, 261.6179, 261.4614, 260.7957, 261.72, 
    261.3616, 260.3889, 260.3169, 255.5694, 256.3455, 256.9419, 256.1194, 
    255.0533, 254.5782, 255.3281, 259.9417, 259.3093, 259.2695, 259.8308, 
    259.5942, 258.7668, 258.626, 258.7383, 258.7349, 258.6116, 258.4587, 
    258.2512, 258.1792, 257.9814, 257.623, 257.2, 256.7036, 256.5117, 
    256.3953, 256.2646, 255.8503, 255.5087, 255.7234, 254.7578, 254.8017, 
    255.141, 255.1878, 255.147, 255.2477, 255.3066, 255.7362, 256.9709, 
    256.248, 256.3706, 256.6252, 256.7004, 257.0854, 257.1113, 257.5481, 
    258.4182, 258.1519, 252.8062, 252.0316, 250.3079, 259.3179, 260.8062, 
    262.3459, 263.0564, 265.627, 268.6943, 250.8284, 253.3797, 250.5906, 
    247.5103, 245.8699, 245.0237, 246.6109, 250.1802, 254.4688, 255.4353, 
    261.0361, 262.311, 264.7292, 267.7578, 270.2922,
  273.8342, 274.5647, 275.2131, 276.0894, 276.8809, 277.0093, 275.301, 
    274.541, 273.4116, 271.0259, 268.6123, 266.8738, 265.5957, 264.6565, 
    263.5845, 262.8835, 262.6292, 262.9651, 262.7542, 258.4424, 262.6802, 
    262.9839, 257.2236, 258.032, 258.1753, 258.6377, 258.3191, 257.6357, 
    256.6958, 256.0972, 256.0164, 256.7581, 256.4478, 255.5482, 255.4961, 
    259.6682, 259.5005, 259.0125, 259.0144, 259.1104, 259.0374, 258.9333, 
    259.0745, 259.6763, 259.5366, 259.2207, 258.958, 258.7739, 258.8616, 
    258.9329, 258.7405, 258.7988, 259.7163, 262.4309, 259.5168, 259.1348, 
    259.4966, 258.7996, 257.9026, 257.9976, 258.2317, 258.5391, 259.844, 
    255.2712, 255.8762, 256.23, 256.4204, 257.1389, 256.6523, 257.3879, 
    258.6973, 255.1522, 255.051, 254.5051, 252.401, 253.6707, 259.6411, 
    259.8293, 261.7161, 264.5452, 268.3042, 271.4277, 250.5556, 256.0188, 
    251.281, 247.1281, 245.9603, 247.1141, 252.0617, 258.1191, 258.7048, 
    262.5015, 264.9153, 267.5181, 270.1975, 272.3882,
  275.8289, 276.562, 277.4153, 278.1787, 278.0679, 278.1919, 266.1104, 
    266.7014, 268.0103, 270.0811, 268.5806, 267.1023, 266.0444, 265.6245, 
    264.4036, 263.5122, 263.1943, 263.5457, 260.79, 259.2715, 259.9045, 
    259.5774, 259.011, 259.9937, 260.2629, 258.7202, 258.3811, 258.5022, 
    258.8521, 258.3677, 257.8782, 257.9187, 258.3008, 258.1467, 257.3301, 
    256.6418, 257.0408, 256.3145, 256.3521, 257.1116, 257.3381, 257.1035, 
    257.6487, 260.9351, 261.2798, 260.875, 260.6846, 260.8928, 261.5884, 
    261.9805, 261.6335, 262.3711, 264.5632, 265.0708, 257.3345, 259.8059, 
    261.4602, 263.2939, 262.2175, 262.2603, 262.8508, 263.106, 263.4482, 
    258.6775, 259.0068, 259.0266, 258.365, 257.6826, 257.019, 258.1665, 
    258.9082, 256.6572, 257.1816, 256.8672, 255.2888, 254.8146, 256.3691, 
    255.9859, 260.4194, 261.7703, 266.4692, 271.4507, 261.9556, 256.9639, 
    253.229, 249.0506, 249.3267, 253.3368, 257.7466, 257.1077, 263.4011, 
    267.0649, 270.5955, 272.8577, 274.6628, 275.3291,
  278.4861, 279.3411, 279.7681, 279.8599, 267.0667, 269.3191, 269.4609, 
    269.4709, 268.5166, 267.9534, 266.9204, 267.4854, 266.6885, 266.7085, 
    263.9043, 263.4624, 262.8755, 262.1924, 261.7295, 261.6172, 261.8389, 
    261.5549, 261.5562, 262.1313, 261.2139, 258.9033, 258.6436, 259.8254, 
    260.7241, 260.0898, 259.1035, 259.106, 259.5427, 259.1663, 257.7524, 
    257.1719, 258.3577, 258.054, 257.8572, 258.4907, 259.0542, 259.0063, 
    258.5649, 258.4011, 258.3027, 258.7236, 258.5435, 258.2715, 258.5261, 
    259.4824, 260.8623, 264.9136, 268.427, 260.9211, 265.7698, 264.6426, 
    262.6296, 263.3318, 263.6287, 263.1553, 263.4116, 263.7288, 263.739, 
    263.4312, 262.28, 261.5718, 260.7649, 260.2952, 259.5544, 258.9543, 
    258.2561, 257.8491, 258.6035, 258.0881, 256.9556, 260.0671, 261.8564, 
    259.5342, 258.1797, 261.8823, 268.3254, 272.1086, 261.8843, 258.2927, 
    254.9096, 252.9612, 255.0587, 258.3735, 268.9607, 268.7444, 270.7788, 
    275.6658, 278.6724, 280.261, 279.896, 278.5269,
  280.7842, 281.1304, 280.9656, 280.6169, 270.5063, 272.1174, 272.7109, 
    270.1309, 270.4734, 270.3823, 269.5906, 268.4912, 267.5081, 267.6653, 
    266.8013, 265.8645, 265.1982, 264.8381, 264.3528, 263.6628, 263.6772, 
    263.6489, 263.9026, 264.2317, 263.9031, 262.9734, 262.0662, 262.041, 
    261.824, 261.2349, 260.1282, 260.728, 261.1753, 261.0588, 260.2627, 
    258.7097, 258.3354, 257.6643, 257.8196, 258.2358, 259.2852, 260.1882, 
    260.2786, 259.7317, 259.4634, 261.5874, 262.4302, 262.4141, 266.4495, 
    267.2993, 267.6768, 269.0339, 270.5967, 263.9922, 267.4663, 267.7588, 
    267.0122, 266.3333, 266.4875, 266.7852, 265.9302, 265.8386, 266.282, 
    266.2317, 266.0693, 264.8259, 263.7192, 262.6445, 261.4751, 260.7434, 
    260.1663, 259.9519, 259.3613, 258.4065, 261.2639, 262.085, 263.2725, 
    260.0188, 259.0996, 264.22, 270.4111, 273.22, 274.8843, 258.5054, 
    260.1504, 256.0225, 274.1357, 273.5627, 273.6143, 276.2271, 280.4268, 
    268.636, 272.5513, 282.1577, 281.8206, 280.9978,
  282.4473, 282.1694, 273.106, 273.3989, 272.3127, 275.5437, 273.2971, 
    272.3921, 272.5669, 271.6763, 270.9438, 270.5164, 269.9026, 269.6377, 
    269.0598, 268.2358, 267.7053, 267.042, 266.5737, 266.3013, 265.9888, 
    265.6458, 265.6956, 265.9846, 266.0247, 265.1155, 264.5879, 264.4578, 
    264.2278, 263.8638, 263.5764, 263.0964, 263.4988, 262.8108, 262.1875, 
    262.1448, 261.3728, 258.7102, 259.3628, 260.1689, 260.9053, 260.9639, 
    260.6814, 260.948, 263.178, 262.97, 262.2566, 262.6169, 268.7546, 
    270.0872, 270.356, 271.7686, 272.8145, 266.8469, 270.6895, 269.4861, 
    268.4187, 267.7566, 266.8591, 267.4609, 267.3274, 266.4741, 266.76, 
    267.6484, 268.0178, 268.2915, 267.6477, 265.9436, 264.4404, 263.5198, 
    262.3582, 261.144, 263.7542, 263.9949, 264.0632, 264.3621, 264.3816, 
    264.7661, 261.5127, 266.5286, 271.1934, 273.8645, 275.501, 258.707, 
    258.0864, 275.2207, 276.5249, 278.0745, 279.1748, 280.418, 282.3315, 
    282.6814, 282.6729, 283.2944, 283.4128, 283.0789,
  282.9053, 282.144, 273.1479, 276.7874, 275.8054, 277.1289, 275.9541, 
    274.0845, 274.3213, 273.6882, 272.4285, 272.0117, 271.4143, 271.1223, 
    270.9836, 270.1104, 269.1245, 269.1458, 268.4458, 267.8464, 267.9697, 
    267.825, 267.3962, 267.4875, 268.0024, 267.2361, 267.5364, 267.1672, 
    266.1997, 266.2483, 265.7817, 265.155, 265.5703, 264.6533, 264.0554, 
    263.7952, 263.1875, 260.8147, 262.103, 262.8848, 263.0249, 262.6995, 
    268.4773, 268.5034, 264.4651, 269.7087, 270.1028, 270.1118, 270.9241, 
    272.0039, 272.3203, 273.4204, 274.3906, 267.3735, 269.7761, 269.1519, 
    268.8279, 269.7012, 268.0337, 267.2344, 268.2925, 268.7812, 269.3042, 
    270.3372, 271.084, 270.8652, 270.5339, 269.437, 267.9487, 266.4426, 
    264.9202, 264.9912, 265.5386, 265.8445, 266.2917, 267.3699, 262.9263, 
    263.3328, 266.301, 266.7717, 270.6047, 274.1067, 275.678, 276.261, 
    276.4521, 277.1492, 278.1702, 279.1233, 279.9995, 280.8376, 281.7874, 
    282.3386, 282.6455, 283.5725, 283.9438, 283.636,
  282.9045, 282.3735, 281.1038, 280.5203, 277.3037, 279.0525, 277.7417, 
    275.3557, 275.6968, 274.4675, 273.5149, 273.4343, 273.5312, 272.54, 
    271.9912, 271.5552, 271.074, 270.8743, 270.5146, 269.9492, 269.6274, 
    269.4114, 269.2776, 269.6782, 270.0605, 270.4749, 270.1624, 269.9761, 
    268.8938, 267.9714, 265.2771, 264.196, 264.6021, 263.9021, 262.3987, 
    263.5691, 263.6953, 262.0403, 266.7314, 268.3408, 268.7444, 269.9463, 
    270.5706, 267.2371, 271.6091, 273.3032, 274.3823, 274.5583, 274.8066, 
    275.1343, 274.9331, 275.4443, 276.0742, 275.8286, 276.0439, 277.0293, 
    278.2095, 278.9468, 279.491, 279.1277, 273.8728, 270.562, 268.2354, 
    270.3579, 272.957, 273.5554, 272.8257, 271.467, 270.1914, 269.2429, 
    268.2373, 268.157, 267.1353, 266.9478, 267.3145, 269.3254, 265.2273, 
    266.4512, 268.2231, 263.7886, 270.0659, 272.9019, 274.741, 276.4075, 
    277.4102, 278.1846, 278.9045, 279.4756, 280.0793, 280.7969, 281.7883, 
    282.8701, 283.3813, 284.1228, 284.3879, 278.7092,
  283.7559, 283.3545, 282.7837, 280.5869, 280.8757, 280.4116, 278.2202, 
    277.239, 276.5259, 275.5293, 275.1367, 275.0164, 274.5686, 274.1621, 
    273.4761, 273.1238, 272.0696, 272.387, 271.7922, 271.948, 271.7432, 
    271.4097, 271.5859, 272.0967, 271.28, 271.616, 271.0508, 271.4404, 
    269.9358, 267.3403, 264.4395, 265.3711, 265.3755, 265.2961, 265.1389, 
    264.4038, 264.9231, 265.9856, 268.385, 271.8984, 273.1367, 273.8127, 
    268.8911, 269.2908, 273.8508, 275.3979, 276.062, 276.29, 276.6399, 
    276.9236, 277.0198, 277.2395, 277.543, 278.0186, 278.468, 279.1013, 
    279.3779, 279.9331, 280.6121, 280.8589, 280.5771, 275.9199, 273.2649, 
    273.0981, 273.0491, 274.2271, 273.9119, 273.0527, 272.011, 271.8599, 
    271.3247, 270.7722, 270.0474, 269.1453, 269.0337, 271.2151, 268.666, 
    269.1479, 268.5591, 267.8899, 269.7661, 273.1802, 274.5044, 276.3457, 
    277.5745, 278.3979, 279.1355, 279.8206, 280.5249, 281.2141, 282.509, 
    283.4661, 284.2432, 284.728, 284.7749, 280.9832,
  282.2061, 284.1316, 281.9365, 281.4346, 281.2065, 280.3269, 279.7422, 
    279.1794, 278.3872, 277.5183, 276.7485, 276.6904, 276.1125, 276.4062, 
    275.6858, 274.6877, 273.9924, 274.2571, 273.658, 273.9897, 274.1716, 
    274.5972, 274.4624, 273.9539, 271.1865, 270.9956, 267.9092, 269.875, 
    271.78, 270.1003, 267.9893, 267.5923, 267.9712, 267.9568, 268.3308, 
    266.8794, 266.5408, 267.2285, 269.7935, 273.5378, 274.5615, 274.8835, 
    269.584, 274.4805, 275.1292, 276.2437, 276.6904, 276.9695, 277.3401, 
    277.6602, 277.949, 278.2776, 278.5686, 278.8621, 279.1499, 279.4299, 
    279.8489, 280.4707, 281.1609, 281.7148, 282.0574, 282.1023, 275.1152, 
    273.6902, 271.8879, 272.0842, 274.5171, 273.9868, 273.4292, 273.5146, 
    273.6118, 272.9182, 272.6682, 271.6421, 271.4771, 272.3616, 270.5156, 
    270.5352, 270.0386, 270.54, 271.7483, 273.1538, 275.1597, 276.3765, 
    277.5918, 278.5825, 279.4712, 280.3308, 281.3215, 281.9346, 282.6389, 
    283.4749, 284.865, 285.3235, 281.7339, 281.979,
  283.3374, 283.231, 282.2725, 281.1487, 280.4971, 279.6936, 280.1855, 
    280.0151, 279.7551, 279.7869, 279.3462, 279.2112, 279.541, 279.7197, 
    279.3936, 277.6807, 276.7996, 277.4438, 276.3367, 275.8672, 274.6187, 
    276.563, 274.8484, 269.3015, 266.3938, 272.2249, 267.6184, 269.5237, 
    271.8721, 271.0146, 270.2854, 270.5103, 269.1562, 269.9192, 270.1453, 
    269.3157, 269.2397, 268.7725, 271.5615, 274.54, 275.4846, 275.5488, 
    275.4246, 275.7151, 276.2085, 276.6943, 277.0066, 277.3193, 277.623, 
    277.917, 278.2488, 278.5769, 278.8911, 279.1978, 279.4958, 279.8774, 
    280.4377, 280.9934, 281.6597, 282.2812, 282.7664, 283.1975, 282.8015, 
    275.0854, 274.8296, 271.7688, 276.2129, 276.26, 275.3469, 274.5569, 
    275.2075, 275.1074, 273.9346, 273.0984, 273.873, 274.6094, 273.2129, 
    273.0068, 273.5708, 273.894, 275.2749, 275.0535, 276.3188, 277.1536, 
    278.1602, 279.2705, 280.0918, 281.0134, 282.3518, 283.2864, 283.7546, 
    284.5874, 285.6216, 286.2051, 285.9155, 285.7007,
  284.2681, 284.092, 280.5999, 276.8193, 279.6501, 282.6411, 281.3286, 
    279.6526, 281.3052, 281.646, 282.4031, 282.8333, 282.8706, 282.5693, 
    282.5713, 281.1118, 280.2422, 280.196, 279.7031, 278.8662, 279.0007, 
    279.2556, 277.3359, 274.0806, 267.5747, 273.5054, 266.3979, 270.0542, 
    272.0183, 270.562, 273.0591, 272.5586, 270.8059, 273.4346, 271.7112, 
    272.8567, 272.1924, 269.7671, 271.2783, 274.3079, 276.0891, 276.3491, 
    276.3716, 276.5859, 276.9106, 277.2192, 277.5598, 277.8638, 278.2356, 
    278.551, 278.8792, 279.2166, 279.5239, 279.8923, 280.2764, 280.6938, 
    281.2214, 281.7393, 282.2856, 282.8635, 283.3997, 283.9937, 283.803, 
    282.4827, 279.5344, 278.5645, 276.1777, 278.4683, 277.5542, 276.7029, 
    276.8418, 276.6826, 276.3508, 279.0659, 274.218, 276.1948, 275.5237, 
    275.7756, 275.9001, 279.1184, 280.1182, 277.3125, 278.1174, 278.7104, 
    279.6648, 281.1477, 281.9399, 282.9287, 284.2979, 285.115, 285.541, 
    285.8794, 286.3818, 287.1318, 287.1926, 287.1143,
  285.7141, 282.1838, 279.6907, 283.1904, 282.9199, 283.0195, 282.7285, 
    282.4797, 284.6028, 285.3301, 286.0806, 283.3638, 285.8049, 285.9158, 
    284.9067, 284.4656, 284.5295, 283.0957, 283.5994, 282.8774, 284.1648, 
    279.4399, 276.6257, 281.1472, 276.6096, 275.5654, 270.2014, 275.7585, 
    276.2722, 276.3508, 275.7361, 273.2454, 274.6211, 275.4644, 273.698, 
    273.9983, 271.5784, 276.457, 274.9578, 274.938, 276.7185, 277.3782, 
    277.4485, 277.6399, 277.9248, 278.3357, 278.7837, 279.1343, 279.5378, 
    279.853, 280.166, 280.4717, 280.741, 281.0984, 281.4453, 281.8545, 
    282.3015, 282.7529, 283.2124, 283.6548, 284.1436, 284.6978, 284.4016, 
    283.3186, 279.334, 277.3367, 274.4919, 276.7002, 278.79, 278.9351, 
    278.791, 279.095, 277.9211, 280.905, 281.3308, 277.9407, 278.5552, 
    277.1492, 278.8433, 280.8608, 281.8945, 280.7629, 280.0181, 281.9756, 
    283.8213, 284.8213, 284.9888, 285.8767, 286.9851, 287.1804, 287.1614, 
    287.2026, 287.5325, 288.05, 287.95, 288.1672,
  282.833, 289.5356, 289.5337, 285.4688, 289.5596, 282.3118, 281.8281, 
    283.9006, 286.8093, 287.4382, 287.9062, 283.3735, 278.634, 286.5701, 
    287.2234, 286.6316, 286.3701, 285.5586, 285.7134, 278.9956, 276.6497, 
    271.3425, 277.2422, 274.4556, 281.4565, 281.2903, 278.5259, 280.1785, 
    278.3347, 278.8735, 277.2065, 274.6079, 277.854, 276.4194, 274.9475, 
    274.3816, 277.916, 279.2878, 276.5676, 276.3689, 277.7463, 278.5576, 
    278.8989, 279.2747, 279.7219, 280.1882, 280.6562, 281.0571, 281.4102, 
    281.7083, 281.9543, 282.2026, 282.427, 282.6848, 282.9727, 283.2883, 
    283.6448, 284.0098, 284.3491, 284.7056, 285.0984, 285.5852, 285.0742, 
    282.2686, 277.9297, 279.8894, 278.4434, 275.7578, 279.1899, 280.6777, 
    281.123, 281.116, 281.0005, 280.979, 281.0994, 280.4387, 280.1238, 
    281.2834, 284.3706, 284.7686, 286.1702, 286.7417, 285.4253, 286.5364, 
    288.0142, 288.1206, 288.085, 288.7827, 289.1077, 288.8047, 288.6123, 
    288.5515, 288.8191, 289.1819, 284.0251, 283.7698,
  286.865, 290.7197, 290.7124, 290.1016, 290.4463, 290.3933, 284.4905, 
    287.5295, 282.6165, 281.5168, 278.3608, 278.4729, 280.6816, 287.0601, 
    290.2227, 288.3301, 287.9885, 287.9507, 284.2917, 277.0242, 271.5544, 
    279.9094, 284.5938, 286.7229, 284.5674, 280.3108, 277.0044, 281.9976, 
    281.8877, 280.8735, 278.2375, 281.0898, 279.8208, 278.4382, 277.1687, 
    280.1758, 281.5588, 282.196, 279.5581, 280.1321, 279.728, 280.5786, 
    281.1631, 281.6604, 282.1323, 282.6089, 283.0198, 283.3774, 283.6685, 
    283.9084, 284.0718, 284.2454, 284.3909, 284.5503, 284.7217, 284.9194, 
    285.1355, 285.3914, 285.6255, 285.8884, 286.1199, 286.2178, 285.2109, 
    285.6614, 280.8459, 278.3831, 280.4575, 278.1003, 278.8853, 283.4539, 
    284.3015, 284.7178, 284.4038, 283.7861, 283.5466, 282.2344, 283.1223, 
    287.9788, 288.8379, 289.9114, 290.5801, 290.7234, 290.3208, 290.4612, 
    290.7622, 290.688, 290.7002, 290.7891, 290.561, 290.1584, 289.8679, 
    289.7051, 289.8198, 289.9827, 287.2705, 285.23,
  289.9604, 291.4575, 291.6235, 291.5254, 291.4685, 291.575, 291.8567, 
    291.0713, 285.0547, 284.3938, 286.3606, 287.4087, 282.1443, 284.249, 
    290.1077, 286.9221, 288.239, 288.8762, 286.5667, 271.1633, 265.2708, 
    281.6714, 283.9944, 273.8684, 267.394, 275.6926, 268.7734, 273.748, 
    280.6492, 281.1047, 280.8894, 285.4795, 284.3679, 283.5234, 279.7126, 
    283.9141, 285.8027, 281.3445, 287.2993, 286.4189, 285.8047, 286.0664, 
    286.2444, 286.3811, 286.5139, 286.5774, 286.5913, 286.6069, 286.582, 
    286.5408, 286.5063, 286.4788, 286.4556, 286.4617, 286.5051, 286.5903, 
    286.7163, 286.8723, 287, 287.1086, 287.1436, 287.0232, 286.8123, 
    287.3293, 282.8179, 281.6965, 281.4377, 281.3257, 280.2922, 286.0757, 
    287.3879, 287.0413, 287.1401, 286.5647, 285.2112, 285.844, 291.5728, 
    292.7739, 293.0027, 292.9021, 292.7432, 292.561, 292.3918, 292.3506, 
    292.3955, 292.3354, 292.2769, 292.0691, 291.6931, 291.2932, 290.9634, 
    290.7876, 290.9695, 291.0881, 290.5728, 287.0825,
  289.248, 289.1667, 289.4365, 292.6047, 292.5093, 292.5288, 292.5977, 
    292.6255, 293.4426, 292.75, 290.0513, 293.4163, 290.0149, 282.6855, 
    285.9114, 290.0864, 288.478, 284.4133, 277.5266, 280.2319, 270.1414, 
    262.3345, 264.5007, 265.3582, 264.7524, 266.6274, 269.9539, 274.1086, 
    279.5659, 283.6418, 284.4187, 286.449, 287.0278, 286.4722, 286.5259, 
    288.3833, 283.7305, 283.0403, 289.9851, 289.802, 289.3447, 289.1602, 
    289.0776, 289.064, 289.0781, 289.0867, 289.071, 289.032, 288.9434, 
    288.8608, 288.7822, 288.6555, 288.4939, 288.3762, 288.2939, 288.2742, 
    288.3069, 288.3596, 288.3633, 288.3125, 288.1934, 288.0142, 287.8687, 
    287.2417, 289.1738, 288.2822, 286.6685, 282.7129, 284.3779, 288.0117, 
    289.8743, 289.7952, 289.6543, 287.9758, 286.6018, 288.0896, 293.6965, 
    294.616, 294.2358, 294.1145, 293.9768, 293.8586, 293.7959, 293.762, 
    293.7297, 293.627, 293.4355, 293.1003, 292.6846, 292.2485, 291.8716, 
    291.6758, 292.0039, 292.3755, 292.8218, 291.7644,
  290.6001, 293.1135, 295.1921, 292.541, 293.2532, 293.2261, 292.9312, 
    292.8545, 293.4902, 292.1465, 290.0754, 293.1453, 296.3967, 289.7349, 
    284.387, 290.3853, 290.1677, 289.2874, 283.4038, 295.1099, 292.0042, 
    268.3818, 264.4038, 267.6741, 269.095, 267.5171, 270.5574, 273.4551, 
    280.9285, 284.1401, 286.325, 287.916, 288.5754, 290.0667, 290.7778, 
    291.842, 292.1626, 291.9062, 292.509, 292.292, 292.0007, 291.6917, 
    291.5088, 291.3479, 291.2227, 291.1272, 291.0688, 290.9824, 290.8674, 
    290.7351, 290.6052, 290.426, 290.2344, 290.085, 289.9695, 289.8792, 
    289.8083, 289.7297, 289.5945, 289.4258, 289.2095, 288.9187, 288.6724, 
    288.7332, 288.8003, 291.7236, 292.2725, 286.7534, 288.2793, 290.3235, 
    291.7041, 292.2981, 291.4387, 290.688, 290.7656, 294.9309, 296.2119, 
    296.0518, 295.5635, 295.366, 295.1895, 295.051, 294.9739, 294.9158, 
    294.8088, 294.6223, 294.3372, 293.9478, 293.5093, 293.082, 292.7427, 
    292.644, 293.2842, 293.4448, 290.9751, 288.1348,
  295.2109, 296.051, 296.0654, 293.7788, 293.7935, 294.4417, 293.7339, 
    293.4954, 294.0745, 292.1028, 291.7729, 293.9099, 296.5627, 297.8889, 
    288.425, 287.4778, 293.9551, 293.3564, 290.6987, 298.615, 299.4165, 
    289.1753, 270.1572, 265.6606, 271.0146, 271.9355, 271.6382, 277.7537, 
    288.5801, 286.4995, 288.7234, 288.9448, 288.8069, 292.5369, 293.6174, 
    294.5823, 294.542, 293.9045, 293.7266, 293.6292, 293.4219, 293.3271, 
    293.2456, 293.1985, 293.1257, 293.0344, 292.9138, 292.7754, 292.6162, 
    292.4336, 292.2344, 292.0217, 291.8171, 291.6321, 291.4475, 291.2649, 
    291.0698, 290.8652, 290.6401, 290.4043, 290.1506, 289.8438, 289.5764, 
    290.0254, 290.5703, 290.3901, 292.8245, 288.8406, 290.3528, 292.2395, 
    293.0454, 293.5098, 292.6985, 292.0386, 292.5449, 296.9434, 296.8594, 
    296.6094, 296.4053, 296.2808, 296.157, 296.0808, 296.0046, 295.8911, 
    295.6877, 295.397, 295.0247, 294.5845, 294.1348, 293.7063, 293.4224, 
    293.3325, 293.9343, 293.7644, 291.4207, 294.5198,
  298.7271, 297.6309, 296.4629, 295.8394, 295.3152, 295.989, 296.3608, 
    295.5266, 295.7795, 296.134, 293.8276, 294.3252, 296.2695, 297.8228, 
    297.7529, 296.2734, 293.5173, 294.364, 297.082, 299.4314, 298.5781, 
    299.8816, 295.95, 285.1477, 282.5657, 288.4475, 283.5234, 281.4404, 
    287.3792, 287.3003, 290.1497, 290.3223, 289.1223, 295.4473, 296.2913, 
    295.8621, 295.4709, 294.9644, 294.864, 294.8616, 294.8855, 294.896, 
    294.8843, 294.8555, 294.7876, 294.6772, 294.5388, 294.3564, 294.1318, 
    293.8965, 293.6428, 293.3757, 293.1177, 292.8523, 292.5906, 292.333, 
    292.0732, 291.804, 291.5293, 291.2603, 290.998, 290.7012, 290.5347, 
    291.0066, 291.8887, 292.626, 294.0718, 290.2083, 289.0906, 293.8169, 
    295.5923, 297.3577, 296.9829, 296.6995, 297.0342, 298.3074, 297.7053, 
    297.4568, 297.332, 297.2432, 297.1411, 297.0354, 296.8694, 296.6392, 
    296.3264, 295.9434, 295.5112, 295.0635, 294.6548, 294.3621, 294.2766, 
    294.575, 295.1885, 293.1423, 296.8391, 297.3726,
  300.7229, 298.021, 294.3838, 295.2778, 296.5796, 296.8257, 296.5657, 
    295.0552, 297.041, 298.4739, 299.5413, 296.0825, 296.7866, 298.4402, 
    301.2144, 301.7112, 299.5139, 298.0098, 295.5886, 298.2803, 298.9368, 
    299.0742, 299.8066, 299.7412, 298.5513, 293.7061, 291.2388, 287.2588, 
    288.7869, 291.1331, 291.2424, 290.5342, 296.9397, 298.4883, 297.6555, 
    296.8379, 296.6238, 296.5164, 296.5488, 296.6355, 296.6831, 296.6575, 
    296.5923, 296.4868, 296.3364, 296.1567, 295.9248, 295.6677, 295.3738, 
    295.0669, 294.7366, 294.4109, 294.0913, 293.7781, 293.4712, 293.1748, 
    292.8796, 292.5781, 292.2891, 292.0308, 291.7869, 291.5498, 291.5562, 
    292.0632, 292.9221, 294.0471, 296.1702, 298.0693, 287.6099, 290.8003, 
    296.6951, 298.9883, 299.033, 299.0488, 298.6672, 299.6514, 298.9553, 
    298.74, 298.4268, 298.2214, 297.989, 297.7505, 297.457, 297.1262, 
    296.7317, 296.3076, 295.8767, 295.4785, 295.2104, 295.0486, 295.0891, 
    295.1599, 295.4116, 296.6697, 299.3088, 300.0852,
  301.3215, 299.0066, 295.7773, 297.8384, 297.8262, 296.291, 297.1265, 
    296.0344, 299.0054, 298.2593, 301.0718, 297.5645, 298.385, 300.8113, 
    302.8352, 301.405, 298.6787, 298.7627, 299.0627, 299.6689, 299.928, 
    299.2773, 298.9304, 299.616, 301.2622, 295.0181, 293.7661, 290.9722, 
    292.4729, 293.8701, 295.2229, 299.0083, 299.2241, 299.396, 298.5852, 
    298.3303, 298.3555, 298.3665, 298.4062, 298.4001, 298.3616, 298.2625, 
    298.1248, 297.9309, 297.7019, 297.4299, 297.1257, 296.792, 296.4514, 
    296.0994, 295.7522, 295.4136, 295.0762, 294.7385, 294.4089, 294.0796, 
    293.762, 293.4573, 293.1606, 292.8809, 292.6382, 292.5071, 292.6763, 
    293.2305, 294.0264, 295.0891, 297.146, 298.572, 293.8376, 288.7485, 
    297.6147, 300.0278, 300.3132, 300.1641, 300.311, 299.905, 300.4517, 
    299.979, 299.2944, 298.9983, 298.6821, 298.3354, 297.9351, 297.5415, 
    297.144, 296.7607, 296.4224, 296.157, 295.9851, 295.8926, 295.9756, 
    296.0525, 297.7922, 299.5784, 300.3164, 301.0742,
  301.8157, 300.1572, 300.0142, 300.5703, 300.2698, 297.4836, 298.3313, 
    298.1831, 299.9958, 299.1377, 299.6921, 298.4568, 298.9292, 301.7781, 
    302.8955, 301.2026, 298.45, 298.707, 299.3911, 299.5347, 298.3662, 
    300.9629, 299.3052, 301.5222, 301.1562, 297.0105, 295.1628, 294.0527, 
    295.0598, 298.6013, 299.855, 300.8047, 300.7322, 300.4658, 300.1255, 
    299.9907, 299.9629, 299.9434, 299.9143, 299.8447, 299.7227, 299.5586, 
    299.354, 299.1035, 298.8027, 298.4792, 298.1389, 297.7825, 297.416, 
    297.043, 296.6702, 296.2998, 295.9175, 295.5413, 295.1746, 294.8354, 
    294.5186, 294.2251, 293.9556, 293.7332, 293.593, 293.6382, 293.9678, 
    294.5818, 295.4155, 296.5901, 298.2578, 299.2051, 296.698, 290.5056, 
    291.4316, 300.8975, 301.749, 300.7202, 301.1692, 302.0918, 301.719, 
    299.8655, 300.0557, 299.6062, 299.3074, 298.9409, 298.5549, 298.1931, 
    297.8203, 297.4644, 297.146, 296.8914, 296.7605, 296.7275, 297.0481, 
    296.8713, 301.4834, 301.3438, 301.2466, 301.8667,
  302.2905, 301.9395, 300.645, 300.9634, 301.98, 302.0859, 299.0632, 
    299.7781, 301.019, 301.166, 300.6636, 303.002, 296.376, 300.0508, 
    299.729, 298.0361, 298.2739, 298.8555, 299.6206, 299.5325, 298.9778, 
    300.9688, 301.4893, 302.0256, 301.5183, 301.0188, 297.1414, 297.3701, 
    297.1653, 300.4663, 301.1296, 301.5601, 301.7014, 301.5544, 301.353, 
    301.1443, 301.0637, 301.0005, 300.9229, 300.783, 300.5942, 300.3616, 
    300.0928, 299.7795, 299.4402, 299.0769, 298.7104, 298.3308, 297.9531, 
    297.5723, 297.209, 296.8433, 296.4888, 296.1533, 295.8518, 295.5964, 
    295.3926, 295.2317, 295.1321, 295.1011, 295.1733, 295.3755, 295.7747, 
    296.3726, 297.1472, 298.1279, 299.3335, 300.2766, 301.0195, 297.9182, 
    293.2622, 298.2898, 302.042, 300.717, 301.0669, 301.3611, 301.2603, 
    300.8594, 300.2363, 300.1301, 299.8035, 299.4058, 299.064, 298.7085, 
    298.3191, 297.97, 297.6943, 297.5088, 297.4558, 297.4954, 297.9158, 
    297.5808, 303.3232, 303.2456, 302.6487, 302.4651,
  302.0625, 301.7119, 301.5068, 301.8655, 302.5537, 301.8584, 298.8652, 
    298.5491, 300.9661, 301.7043, 299.4199, 302.0867, 294.0217, 299.3127, 
    298.5256, 299.4746, 299.4724, 299.6836, 300.1887, 299.9851, 299.2617, 
    302.3757, 301.9475, 301.4412, 301.2766, 300.916, 300.6406, 298.8137, 
    299.1575, 297.8652, 301.6819, 301.9863, 299.8379, 302.136, 301.9121, 
    301.8059, 301.667, 301.5564, 301.3948, 301.1802, 300.9214, 300.6326, 
    300.3203, 299.9883, 299.6477, 299.3052, 298.9731, 298.6453, 298.3296, 
    298.0352, 297.7573, 297.4983, 297.2637, 297.0642, 296.8997, 296.7791, 
    296.7146, 296.7102, 296.7676, 296.9023, 297.1348, 297.4487, 297.8477, 
    298.3621, 298.9556, 299.6064, 300.3037, 300.8896, 301.3049, 301.4792, 
    301.325, 301.2517, 297.4954, 298.2905, 300.7407, 300.9167, 300.6272, 
    300.645, 300.6267, 300.5503, 300.343, 299.8867, 299.4612, 299.1104, 
    298.7639, 298.4524, 298.2288, 298.1016, 298.0989, 298.1985, 298.614, 
    298.3652, 303.1699, 303.4927, 302.46, 302.4045,
  300.8191, 300.7375, 299.4463, 301.1021, 302.7871, 300.5901, 298.4011, 
    299.3362, 300.5417, 301.2588, 293.1731, 300.114, 299.7131, 299.668, 
    300.3059, 300.303, 299.9949, 300.1567, 300.6289, 300.9636, 301.3696, 
    300.2261, 301.9106, 301.6875, 301.4023, 301.1321, 301.0903, 299.9915, 
    300.6829, 298.6626, 301.8582, 302.1821, 302.637, 300.9429, 302.0789, 
    301.9187, 301.8015, 301.6492, 301.468, 301.2393, 301.0029, 300.7385, 
    300.4795, 300.2024, 299.9341, 299.6667, 299.4219, 299.1929, 298.9873, 
    298.8015, 298.6401, 298.5007, 298.3916, 298.3052, 298.248, 298.219, 
    298.2288, 298.2798, 298.3816, 298.5405, 298.7722, 299.0681, 299.4136, 
    299.8093, 300.2227, 300.6025, 300.9241, 301.1567, 301.2917, 301.3706, 
    301.4763, 301.9033, 302.7356, 300.6089, 300.5186, 299.2864, 298.0637, 
    297.4082, 298.1758, 299.8152, 300.5322, 300.4102, 299.9717, 299.5762, 
    299.27, 299.0239, 298.8538, 298.7891, 298.8071, 298.936, 299.2854, 
    299.3186, 301.4558, 299.9595, 300.2578, 300.7917,
  299.8682, 299.1863, 297.3433, 299.4663, 300.8157, 300.5452, 299.5688, 
    299.9653, 301.3098, 298.2014, 290.3813, 296.3184, 299.9521, 299.314, 
    300.0244, 300.3979, 300.4749, 300.7278, 301.0305, 301.3423, 301.7776, 
    302.1975, 301.8459, 301.6819, 301.53, 301.4968, 301.6089, 300.6619, 
    301.1426, 301.9331, 301.9741, 302.4634, 302.8748, 300.8354, 302.1777, 
    302.03, 301.9385, 301.7974, 301.6514, 301.4854, 301.3276, 301.1602, 
    300.9954, 300.8228, 300.6538, 300.4924, 300.343, 300.2092, 300.0908, 
    299.9907, 299.9016, 299.8303, 299.7676, 299.7183, 299.6843, 299.6721, 
    299.676, 299.7041, 299.7612, 299.8589, 299.9868, 300.1509, 300.3306, 
    300.5308, 300.7488, 300.9558, 301.1025, 301.1804, 301.229, 301.3066, 
    301.481, 301.7664, 302.0747, 302.0886, 298.2153, 301.3462, 301.719, 
    301.2109, 301.395, 301.6411, 300.3484, 300.5457, 300.45, 300.1418, 
    299.8203, 299.6843, 299.5706, 299.5383, 299.5667, 299.6602, 299.8855, 
    300.1497, 300.9355, 297.825, 298.687, 299.5344,
  299.1877, 299.0815, 299.0537, 296.9553, 297.5037, 300.0662, 297.4927, 
    298.6841, 301.7039, 298.5146, 290.2134, 295.1816, 299.822, 298.1406, 
    300.6479, 300.9702, 301.1733, 301.3481, 301.5022, 301.6729, 301.6628, 
    301.7942, 301.3967, 301.5876, 301.6924, 301.8127, 301.9121, 302.2278, 
    302.2634, 302.2185, 302.3774, 303.0186, 302.9614, 299.1941, 302.3511, 
    302.252, 302.1943, 302.0811, 301.98, 301.873, 301.7803, 301.686, 
    301.5942, 301.5005, 301.407, 301.311, 301.2246, 301.1377, 301.0576, 
    300.9783, 300.9092, 300.843, 300.7812, 300.7222, 300.6733, 300.627, 
    300.5903, 300.5613, 300.5481, 300.5466, 300.5596, 300.5925, 300.6455, 
    300.7129, 300.8015, 300.8887, 300.9595, 301.0022, 301.0562, 301.1406, 
    301.2673, 301.3972, 301.4246, 301.5054, 301.594, 299.9475, 297.6687, 
    297.0786, 302.7307, 301.1504, 301.1458, 300.4182, 300.6924, 300.7971, 
    300.3943, 300.3308, 300.2742, 300.2468, 300.2744, 300.3677, 300.5618, 
    300.8555, 301.0667, 298.8977, 298.4348, 299.4658,
  301.4866, 301.6533, 299.6008, 296.916, 297.28, 298.6475, 298.4104, 
    297.5205, 298.6746, 298.019, 293.9124, 300.2354, 301.5723, 301.292, 
    301.1316, 301.3052, 301.4692, 301.637, 301.7629, 301.8521, 301.8137, 
    301.7219, 301.6526, 301.7649, 301.8909, 302.0742, 302.2673, 299.3247, 
    302.6724, 302.4739, 302.9714, 299.0056, 302.9109, 302.5764, 302.3186, 
    302.4231, 302.3945, 302.2744, 302.1807, 302.0872, 302.0249, 301.9578, 
    301.8811, 301.7996, 301.7136, 301.6216, 301.5176, 301.4072, 301.2815, 
    301.1584, 301.0398, 300.9358, 300.843, 300.7627, 300.687, 300.6187, 
    300.5588, 300.5137, 300.479, 300.4351, 300.3855, 300.3687, 300.3853, 
    300.4314, 300.4915, 300.5371, 300.5815, 300.6375, 300.7058, 300.79, 
    300.8855, 300.9758, 301.0146, 301.0264, 301.156, 301.4102, 292.27, 
    298.9817, 299.5093, 297.9905, 298.8889, 301.2014, 300.396, 300.7844, 
    300.7659, 300.7446, 300.7256, 300.7271, 300.7151, 300.77, 300.855, 
    300.9824, 300.9846, 301.2563, 299.2747, 299.8752,
  301.3027, 301.4868, 301.4248, 298.0159, 298.1887, 299.2104, 299.2275, 
    298.2493, 295.5518, 294.646, 300.8127, 301.7, 301.9473, 301.2012, 
    301.2869, 301.5164, 301.6301, 301.7144, 301.7756, 301.8118, 301.8147, 
    301.7847, 301.8149, 301.8987, 302.0249, 302.1797, 302.3826, 300.9399, 
    302.6316, 302.5415, 300.3904, 298.1838, 302.7297, 302.5281, 302.5164, 
    302.5237, 302.395, 302.2449, 302.1382, 302.0029, 301.8657, 301.6978, 
    301.5151, 301.3225, 301.1267, 300.9199, 300.7097, 300.4978, 300.2969, 
    300.1199, 299.95, 299.8032, 299.6702, 299.5425, 299.4084, 299.2905, 
    299.2, 299.1194, 299.0713, 299.0366, 299.0085, 298.9878, 298.9946, 
    299.0605, 299.1646, 299.2903, 299.4243, 299.5803, 299.7649, 299.9763, 
    300.1965, 300.376, 300.5142, 300.6357, 300.7649, 300.8928, 294.6042, 
    299.8789, 300.5576, 298.646, 302.9595, 302.011, 300.4136, 300.5684, 
    300.5305, 300.6101, 300.5808, 300.6455, 300.594, 300.5891, 300.6079, 
    300.7021, 300.7473, 300.8142, 300.9202, 301.0869,
  301.1421, 301.3474, 301.3242, 298.9619, 298.6035, 299.4453, 299.4719, 
    298.0061, 294.0273, 293.9424, 296.1042, 301.5793, 301.2344, 300.9573, 
    301.3271, 301.449, 301.501, 301.5769, 301.6555, 301.7234, 301.7805, 
    301.8325, 301.9016, 301.979, 302.0793, 302.2004, 302.3345, 300.0847, 
    302.8369, 302.6685, 299.4006, 300.2061, 303.0215, 302.5774, 302.6216, 
    302.6492, 302.5593, 302.4082, 301.8848, 301.5151, 301.2805, 300.9927, 
    300.7334, 300.4729, 300.2273, 299.9863, 299.7551, 299.5356, 299.3262, 
    299.1206, 298.9192, 298.7197, 298.5332, 298.3501, 298.1616, 297.9868, 
    297.8203, 297.6597, 297.4819, 297.302, 297.1069, 296.9351, 296.7388, 
    296.6277, 296.5457, 296.573, 296.6748, 296.8591, 297.1709, 297.7209, 
    298.4255, 299.135, 299.6614, 300.0244, 300.0371, 294.2273, 299.3135, 
    300.4651, 300.8289, 300.6628, 301.5408, 303.4136, 301.8762, 300.5698, 
    300.3909, 300.0859, 299.842, 299.9443, 299.8328, 299.7925, 299.7876, 
    299.9368, 300.0725, 300.2729, 300.5217, 300.8501,
  300.8689, 301.2317, 301.4858, 299.1394, 298.1328, 299.5894, 298.8154, 
    297.2883, 291.9937, 295.2883, 296.5859, 300.5679, 300.9685, 301.1443, 
    301.3132, 301.3489, 301.3704, 301.4045, 301.4358, 301.4646, 301.5007, 
    301.5515, 301.6245, 301.7227, 301.8604, 302.0413, 302.2236, 299.7627, 
    301.3989, 302.6929, 301.2004, 301.4084, 297.5505, 302.7358, 302.5198, 
    302.6243, 302.9893, 299.9783, 302.2825, 301.8596, 301.6411, 301.5039, 
    301.3284, 301.1641, 301.0088, 300.8464, 300.687, 300.5281, 300.3801, 
    300.2234, 300.0664, 299.9041, 299.7454, 299.5969, 299.4514, 299.3054, 
    299.1624, 299.0247, 298.8635, 298.7014, 298.543, 298.3889, 298.2412, 
    298.137, 298.0676, 298.0715, 298.0864, 298.1414, 298.2312, 298.4521, 
    298.7178, 299.1191, 299.5076, 299.6677, 299.075, 294.8621, 300.2119, 
    301.0842, 301.3691, 301.7595, 301.5117, 302.3347, 302.8713, 301.3113, 
    300.8079, 300.8098, 300.3442, 299.7339, 299.8811, 299.7646, 299.741, 
    299.8081, 299.8765, 300.0298, 300.2219, 300.5386,
  300.4453, 300.96, 301.334, 300.9851, 298.5132, 298.5278, 298.3174, 297.561, 
    294.9031, 294.6829, 294.9368, 300.6333, 301.0847, 301.1438, 301.1665, 
    301.1711, 301.1572, 301.1721, 301.1882, 301.2012, 301.2239, 301.272, 
    301.3567, 301.479, 301.646, 301.8252, 302.0024, 302.4048, 300.0908, 
    302.5857, 302.4814, 302.3823, 302.3992, 302.4971, 302.4082, 302.4392, 
    302.4675, 298.2092, 295.9429, 302.0645, 302.0391, 302.1262, 302.0835, 
    302.0166, 301.9683, 301.8948, 301.8164, 301.741, 301.6611, 301.5728, 
    301.479, 301.3916, 301.2969, 301.1946, 301.0872, 300.9663, 300.8218, 
    300.6553, 300.4641, 300.2622, 300.0542, 299.853, 299.6697, 299.519, 
    299.3853, 299.2783, 299.1792, 299.1077, 299.0801, 299.0991, 299.1428, 
    299.3018, 299.6006, 299.7646, 298.6965, 294.2991, 300.4241, 301.0742, 
    301.5586, 302.0022, 302.0264, 301.7664, 301.1228, 300.8049, 300.9541, 
    300.5308, 301.7512, 299.6731, 299.9497, 299.8135, 299.7292, 299.665, 
    299.6367, 299.6648, 299.7803, 300.0354,
  299.5593, 300.2129, 300.7014, 299.9243, 297.7815, 296.614, 296.5681, 
    297.0808, 295.4858, 294.4976, 297.29, 300.6106, 300.8091, 300.7341, 
    300.7, 300.7009, 300.6477, 300.6538, 300.6677, 300.6917, 300.7395, 
    300.8291, 300.9609, 301.1436, 301.3767, 301.5898, 301.7229, 301.8691, 
    302.1733, 302.3286, 302.3433, 302.3838, 302.4924, 302.2686, 302.2217, 
    302.2129, 302.0615, 301.7239, 300.6272, 296.7664, 301.8088, 302.0823, 
    302.0947, 302.1011, 302.1023, 302.0908, 302.0774, 302.0547, 302.0352, 
    302.0037, 301.9661, 301.9172, 301.8562, 301.7659, 301.6536, 301.5093, 
    301.3306, 301.1145, 300.8667, 300.5928, 300.3105, 300.0178, 299.7175, 
    299.4231, 299.1487, 298.9058, 298.7014, 298.5417, 298.4263, 298.3811, 
    298.4226, 298.6299, 299.0066, 299.4756, 298.759, 291.6177, 298.2451, 
    300.5029, 301.1597, 301.7949, 301.739, 300.6272, 300.2791, 299.9541, 
    300.1868, 300.8906, 299.2366, 298.8955, 299.4873, 299.1616, 298.9714, 
    298.8098, 298.7268, 298.709, 298.8242, 299.0918,
  298.5574, 299.2708, 299.9185, 299.1382, 298.1201, 295.4553, 295.9612, 
    295.457, 295.0403, 293.6235, 296.6772, 300.4241, 300.4805, 300.2112, 
    300.1147, 300.1594, 300.0364, 300.0303, 300.0254, 300.05, 300.1157, 
    300.2415, 300.4146, 300.6348, 300.8958, 301.1646, 301.3862, 301.551, 
    301.7512, 301.8669, 301.9778, 302.0596, 302.0842, 302.0034, 301.9719, 
    301.9539, 301.8643, 301.2227, 301.3953, 301.1826, 301.5659, 301.6917, 
    301.688, 301.7114, 301.7305, 301.7546, 301.7742, 301.7903, 301.8074, 
    301.822, 301.833, 301.8323, 301.8203, 301.7759, 301.6904, 301.5554, 
    301.3599, 301.1064, 300.7971, 300.4436, 300.0581, 299.6499, 299.2251, 
    298.8083, 298.4229, 298.0732, 297.771, 297.5264, 297.3516, 297.2805, 
    297.3364, 297.5706, 297.9783, 298.6067, 298.6848, 297.6924, 291.7578, 
    299.5654, 300.4695, 300.3684, 300.4646, 299.8157, 299.6626, 299.95, 
    298.5608, 298.7666, 298.771, 298.98, 298.7671, 298.3938, 298.1055, 
    297.8684, 297.741, 297.6997, 297.812, 298.0815,
  297.5339, 298.2754, 299.1863, 298.8708, 294.3159, 294.3899, 295.5127, 
    295.0791, 294.9319, 295.5237, 296.0503, 300.5012, 300.7229, 300.0039, 
    299.6208, 299.7288, 299.5088, 299.4109, 299.3391, 299.3159, 299.3306, 
    299.4011, 299.5093, 299.6648, 299.8496, 300.0596, 300.2769, 300.511, 
    300.8113, 301.116, 301.4348, 301.6997, 301.8679, 301.9937, 302.1084, 
    302.2271, 300.3115, 301.1399, 301.0081, 300.821, 301.1697, 301.0996, 
    301.0977, 301.1421, 301.1914, 301.2339, 301.2705, 301.2917, 301.3215, 
    301.3577, 301.4004, 301.4238, 301.4399, 301.4395, 301.4126, 301.3242, 
    301.1533, 300.8972, 300.5569, 300.1416, 299.6748, 299.1672, 298.6406, 
    298.1223, 297.6394, 297.1914, 296.8059, 296.4915, 296.2456, 296.103, 
    296.0806, 296.2175, 296.5574, 297.2209, 298.1462, 297.6829, 286.0315, 
    291.4402, 299.1558, 299.2815, 298.8997, 299.1318, 299.3679, 298.5535, 
    296.9407, 295.8125, 298.0139, 298.7012, 298.2246, 297.717, 297.3379, 
    297.0376, 296.8464, 296.7622, 296.8389, 297.071,
  296.3694, 297.0513, 298.0693, 297.9155, 293.863, 294.8218, 296.2466, 
    295.624, 296.6414, 296.4185, 296.2925, 300.6392, 301.6597, 297.8508, 
    299.0366, 299.3723, 299.0259, 298.7817, 298.5906, 298.4307, 298.323, 
    298.2761, 298.2722, 298.3445, 298.4626, 298.6265, 298.8616, 299.2017, 
    299.6548, 300.1636, 300.7266, 301.2666, 301.7207, 302.3777, 300.2849, 
    300.9102, 301.1067, 301.6453, 300.0688, 300.0605, 300.2161, 300.3398, 
    300.3511, 300.3975, 300.446, 300.4937, 300.5168, 300.5315, 300.5435, 
    300.5801, 300.6194, 300.6523, 300.6755, 300.6963, 300.7012, 300.6643, 
    300.5454, 300.3401, 300.03, 299.6328, 299.1624, 298.6357, 298.0791, 
    297.5161, 296.9561, 296.4109, 295.915, 295.4868, 295.1155, 294.8584, 
    294.7119, 294.7192, 294.9072, 295.302, 296.2324, 295.957, 292.8875, 
    278.6538, 292.1614, 298.7129, 297.9448, 298.4912, 297.7278, 295.5869, 
    296.272, 294.9734, 298.1565, 298.3027, 297.6067, 297.1033, 296.6619, 
    296.2981, 296.0183, 295.8611, 295.8457, 295.9966,
  295.2034, 295.759, 296.7336, 296.3992, 294.6289, 296.051, 296.1362, 
    296.3521, 294.2349, 296.3918, 299.4429, 300.8149, 301.6106, 297.1016, 
    298.7388, 299.0417, 298.6086, 298.2441, 297.9207, 297.6079, 297.3452, 
    297.135, 296.9902, 296.9517, 297.0005, 297.1392, 297.4126, 297.8423, 
    298.4282, 299.1296, 299.9385, 300.7373, 301.3765, 300.155, 298.7625, 
    300.1047, 300.1721, 301.1179, 299.8323, 299.5691, 299.3008, 299.4377, 
    299.4895, 299.5054, 299.5071, 299.5125, 299.4966, 299.4797, 299.4585, 
    299.4526, 299.4604, 299.4709, 299.4924, 299.5293, 299.5725, 299.593, 
    299.5742, 299.5103, 299.3645, 299.1301, 298.8035, 298.3831, 297.9075, 
    297.3945, 296.8447, 296.2603, 295.6675, 295.1011, 294.5891, 294.1746, 
    293.8816, 293.709, 293.738, 293.9573, 294.5083, 294.1426, 292.4036, 
    291.2566, 280.8931, 294.4268, 298.1628, 299.3591, 295.8743, 295.0056, 
    294.7129, 294.4646, 297.7295, 297.6516, 297.0735, 296.583, 296.0925, 
    295.6682, 295.3047, 295.0542, 294.9119, 294.9436,
  294.1904, 294.5852, 295.3713, 294.9639, 294.7678, 294.3208, 296.0366, 
    295.5854, 293.623, 297.0283, 300.5598, 300.7249, 301.395, 296.4304, 
    298.5618, 298.647, 298.2051, 297.7937, 297.4155, 297.0413, 296.6702, 
    296.3264, 296.0244, 295.8413, 295.7737, 295.8208, 296.0347, 296.4387, 
    297.0862, 297.9543, 299.0161, 300.1646, 300.2686, 299.8362, 298.9407, 
    298.2949, 298.4883, 298.7979, 298.8284, 295.9495, 298.9871, 298.5972, 
    298.5522, 298.5454, 298.4915, 298.4514, 298.3894, 298.3242, 298.2493, 
    298.1824, 298.1333, 298.1038, 298.0854, 298.1003, 298.1418, 298.2039, 
    298.2546, 298.3186, 298.3518, 298.323, 298.2205, 298.0127, 297.7075, 
    297.3113, 296.8586, 296.3569, 295.8123, 295.2219, 294.6196, 294.0532, 
    293.5698, 293.1738, 292.9299, 292.9072, 293.3198, 294.1741, 294.585, 
    293.2773, 278.6538, 291.0432, 296.8918, 298.1204, 296.6641, 295.2471, 
    292.2307, 294.6235, 297.5378, 297.0789, 296.6199, 296.1677, 295.6978, 
    295.2522, 294.842, 294.5017, 294.2156, 294.0811,
  293.3872, 293.5203, 294.0957, 293.7258, 296.0208, 291.6846, 293.9514, 
    293.9685, 295.7886, 297.3718, 300.0938, 300.2937, 294.082, 298.9478, 
    298.5522, 298.2036, 297.7278, 297.2622, 296.8315, 296.4368, 296.0518, 
    295.6675, 295.2832, 294.9709, 294.7363, 294.6453, 294.7473, 295.041, 
    295.6917, 296.7, 297.8132, 296.0776, 296.3823, 298.1125, 297.6443, 
    294.9265, 295.334, 297.5007, 297.5273, 296.6138, 296.5579, 297.76, 
    297.4917, 297.5479, 297.4788, 297.418, 297.3367, 297.2368, 297.1272, 
    297.0024, 296.8845, 296.7935, 296.7288, 296.6855, 296.675, 296.7107, 
    296.7852, 296.8835, 296.9983, 297.1069, 297.1926, 297.2046, 297.1172, 
    296.9109, 296.5981, 296.1948, 295.7319, 295.2112, 294.6301, 294.0222, 
    293.4358, 292.8855, 292.427, 292.1196, 292.0776, 292.6414, 293.5186, 
    292.5112, 277.7905, 291.5474, 295.7622, 296.0469, 295.7559, 293.3914, 
    291.51, 297.2976, 296.9636, 296.5544, 296.1367, 295.7561, 295.3557, 
    294.9575, 294.5708, 294.187, 293.8176, 293.5317,
  292.8875, 292.7424, 293.0535, 292.3894, 292.3374, 291.749, 292.9165, 
    291.4246, 290.7771, 296.7434, 299.2544, 299.3867, 297.0752, 298.4631, 
    297.7854, 297.4822, 297.0593, 296.5913, 296.136, 295.7021, 295.2947, 
    294.8977, 294.4802, 294.1213, 293.8232, 293.6038, 293.5652, 293.7278, 
    294.2979, 295.2925, 296.5469, 294.8489, 293.7183, 294.5442, 294.5801, 
    292.8506, 294.9976, 296.8416, 296.1001, 293.8535, 293.2007, 296.8782, 
    296.3782, 296.4387, 296.373, 296.3467, 296.2825, 296.197, 296.0884, 
    295.9563, 295.7979, 295.6436, 295.5122, 295.415, 295.3542, 295.3391, 
    295.3713, 295.4424, 295.5515, 295.6951, 295.843, 295.9802, 296.0574, 
    296.0435, 295.9238, 295.6782, 295.3269, 294.8879, 294.3748, 293.8027, 
    293.1919, 292.5645, 292.0049, 291.574, 291.3608, 291.7832, 292.5876, 
    291.9041, 276.1228, 292.7778, 295.2786, 295.5991, 292.3242, 292.0798, 
    296.7512, 296.6804, 296.1687, 295.8252, 295.5112, 295.1868, 294.8403, 
    294.4946, 294.1562, 293.8052, 293.458, 293.1479,
  292.3274, 292.1521, 292.2812, 292.1274, 289.8801, 291.1545, 290.7493, 
    288.5317, 287.5342, 298.4307, 298.3267, 298.1509, 297.8164, 297.0337, 
    296.6052, 296.325, 295.9707, 295.561, 295.0964, 294.6365, 294.2671, 
    293.8772, 293.4426, 293.0669, 292.7739, 292.585, 292.5105, 292.5293, 
    292.9172, 293.8308, 295.0696, 293.1904, 291.9053, 291.7542, 292.4204, 
    291.4824, 293.8574, 295.3457, 294.304, 293.4067, 291.3872, 295.9526, 
    295.2571, 295.2163, 295.123, 295.1025, 295.0762, 295.0168, 294.9351, 
    294.8086, 294.6399, 294.4519, 294.2812, 294.1296, 294.0161, 293.9604, 
    293.9595, 294.0029, 294.0842, 294.2107, 294.3567, 294.5234, 294.6792, 
    294.8015, 294.8413, 294.7646, 294.5637, 294.2444, 293.8313, 293.3328, 
    292.7578, 292.1172, 291.5029, 290.9814, 290.6411, 291.0134, 291.52, 
    291.6206, 278.4736, 292.0403, 294.3132, 294.5059, 290.4988, 290.9448, 
    295.7759, 295.3684, 294.9556, 294.7134, 294.5208, 294.3123, 294.0686, 
    293.7837, 293.5007, 293.1851, 292.8704, 292.5708,
  291.5715, 291.4182, 291.5383, 292.1353, 291.1467, 291.0496, 288.8518, 
    286.0676, 287.7117, 297.667, 296.2329, 295.9124, 295.5125, 295.1506, 
    294.9834, 294.791, 294.5505, 294.2776, 293.9216, 293.5042, 293.2041, 
    292.8691, 292.4019, 291.9492, 291.5732, 291.3196, 291.2002, 291.2017, 
    291.457, 292.145, 293.3853, 291.7578, 290.3086, 290.0676, 289.7903, 
    290.8203, 292.0017, 293.0229, 292.6357, 292.9741, 289.2739, 295.1865, 
    294.3408, 294.2056, 294.0825, 293.9983, 293.9211, 293.876, 293.8201, 
    293.6729, 293.4675, 293.2485, 293.0276, 292.8203, 292.6492, 292.5439, 
    292.4907, 292.4927, 292.5461, 292.6433, 292.7627, 292.927, 293.1047, 
    293.2876, 293.4233, 293.4753, 293.4226, 293.2463, 292.968, 292.6008, 
    292.1223, 291.5376, 290.9189, 290.4121, 290.03, 290.0918, 289.1763, 
    284.8862, 286.8066, 291.5244, 293.5977, 292.5718, 291.0852, 294.3865, 
    294.5225, 293.7959, 293.4736, 293.2842, 293.1216, 293.0049, 292.8596, 
    292.6663, 292.4729, 292.2593, 292.0229, 291.802,
  290.626, 290.5706, 290.5889, 290.8362, 290.1946, 289.0696, 285.6631, 
    286.4639, 295.9551, 296.053, 294.7803, 294.1067, 293.7656, 293.5457, 
    293.3811, 293.1709, 292.9763, 292.7756, 292.5479, 292.2051, 291.9102, 
    291.6467, 291.2285, 290.8003, 290.4268, 290.0845, 289.8403, 289.7603, 
    289.9263, 290.5247, 291.7656, 289.5474, 288.5249, 288.7124, 290.8975, 
    291.1514, 289.8264, 290.3618, 291.4509, 290.4104, 287.614, 294.2449, 
    293.5535, 293.3445, 293.1729, 293.0828, 293.0522, 292.9927, 292.7991, 
    292.6323, 292.387, 292.1208, 291.8564, 291.6035, 291.3796, 291.2056, 
    291.094, 291.0295, 291.0237, 291.0706, 291.1418, 291.2708, 291.4155, 
    291.584, 291.7446, 291.8633, 291.9102, 291.8718, 291.7241, 291.4888, 
    291.146, 290.7043, 290.1636, 289.614, 289.239, 289.585, 287.6665, 
    284.4482, 287.9141, 289.5083, 292.7727, 290.8889, 290.8589, 293.21, 
    292.5637, 292.1409, 291.9041, 291.7017, 291.5378, 291.4487, 291.3623, 
    291.2461, 291.1213, 290.9875, 290.8528, 290.7278,
  289.657, 289.7864, 290.0081, 290.5852, 290.813, 290.9639, 292.0957, 
    293.7847, 294.7703, 295.0295, 294.0928, 293.2561, 292.6838, 292.3352, 
    292.1194, 291.8855, 291.6763, 291.4033, 291.1777, 290.9761, 290.7241, 
    290.2996, 289.9441, 289.5359, 289.1672, 288.8171, 288.5684, 288.45, 
    288.4939, 288.9546, 289.6409, 289.2725, 289.5139, 289.6421, 289.5676, 
    289.8452, 290.1555, 289.1326, 289.8699, 289.0828, 286.0964, 293.6841, 
    292.8921, 292.4084, 292.0693, 291.8845, 291.8665, 292.0823, 291.7698, 
    291.5752, 291.2803, 290.9685, 290.6587, 290.3682, 290.114, 289.8906, 
    289.7122, 289.5708, 289.4836, 289.4692, 289.491, 289.5503, 289.6304, 
    289.7429, 289.8792, 290.0042, 290.0791, 290.1135, 290.0706, 289.9419, 
    289.731, 289.4399, 289.0315, 288.5774, 288.1353, 288.5867, 287.553, 
    283.3235, 286.4844, 290.4089, 290.6108, 290.0244, 291.6589, 291.7922, 
    290.9587, 290.5505, 290.2686, 290.0342, 289.8721, 289.8118, 289.7637, 
    289.6794, 289.5786, 289.5076, 289.4607, 289.4585,
  287.8772, 288.0171, 288.1597, 288.5776, 289.3079, 290.2744, 291.302, 
    291.9229, 292.6172, 291.6917, 291.4316, 291.5203, 291.4153, 291.3362, 
    291.1782, 290.7649, 290.3474, 290.2146, 290.1521, 289.9585, 289.7944, 
    289.2141, 288.8296, 288.4487, 288.0515, 287.6453, 287.3215, 287.1162, 
    287.0239, 287.0947, 287.2458, 287.3428, 287.551, 287.6809, 287.7473, 
    287.9661, 288.3206, 288.9182, 286.9036, 285.5938, 290.9834, 292.4324, 
    291.7456, 291.053, 290.5901, 290.4167, 290.6396, 291.075, 291.1829, 
    290.6086, 290.1863, 289.7876, 289.437, 289.1106, 288.8291, 288.5542, 
    288.3389, 288.1304, 287.9766, 287.8826, 287.8374, 287.8137, 287.8296, 
    287.8745, 287.9519, 288.0276, 288.084, 288.1309, 288.1604, 288.1077, 
    287.9827, 287.8062, 287.5386, 287.2886, 286.967, 287.3276, 287.0281, 
    281.3774, 286.1357, 288.5059, 288.1355, 289.8823, 290.4285, 289.8821, 
    289.366, 289.0454, 288.7839, 288.5935, 288.4419, 288.3777, 288.2307, 
    288.113, 287.9744, 287.8184, 287.7996, 287.7278,
  285.7881, 285.7339, 285.624, 285.5945, 285.7371, 286.1641, 286.7119, 
    286.4016, 286.3137, 285.6648, 285.7834, 286.8547, 287.4827, 287.8625, 
    288.1545, 287.636, 286.9883, 286.9951, 287.4309, 287.5403, 288.0967, 
    287.7461, 287.386, 287.0554, 286.7559, 286.5051, 286.271, 286.0161, 
    285.8098, 285.6372, 285.5654, 285.5713, 285.6602, 285.7544, 285.8818, 
    286.0583, 286.3508, 286.907, 287.4934, 287.9773, 289.2944, 288.7061, 
    289.1792, 289.0283, 288.9324, 289.2131, 289.7222, 284.8342, 290.5811, 
    289.7776, 289.1804, 288.6475, 288.2334, 287.8838, 287.5867, 287.2947, 
    287.0449, 286.7915, 286.5894, 286.4277, 286.3281, 286.2239, 286.1497, 
    286.1318, 286.134, 286.1426, 286.1567, 286.1846, 286.2385, 286.2327, 
    286.1638, 286.074, 285.895, 285.7952, 285.6077, 285.8853, 285.8748, 
    280.2847, 284.4243, 287.2046, 286.8262, 287.7209, 289.0242, 287.7124, 
    287.165, 286.772, 286.4951, 286.3945, 286.4377, 286.6875, 286.8872, 
    286.7649, 286.4414, 286.3997, 286.1414, 285.9255,
  283.9133, 283.709, 283.4951, 283.3713, 283.2874, 283.2971, 283.4697, 
    283.3638, 283.4399, 283.1101, 282.9414, 283.9211, 284.3804, 284.4546, 
    284.2642, 283.9724, 283.7656, 283.6543, 284.0088, 284.1594, 285.4692, 
    285.5811, 285.4873, 285.2512, 285.0012, 284.7671, 284.7017, 284.5984, 
    284.509, 284.436, 284.3931, 284.3328, 284.3345, 284.3518, 284.3923, 
    284.5522, 284.8779, 285.4932, 286.123, 286.8176, 287.9983, 287.2009, 
    287.55, 287.3606, 287.5759, 287.8733, 281.9199, 289.1057, 289.5178, 
    288.8479, 288.1572, 287.6213, 287.2356, 286.8428, 286.4009, 286.0557, 
    285.7646, 285.4893, 285.2686, 285.0942, 284.9651, 284.8313, 284.6831, 
    284.6077, 284.5605, 284.4888, 284.467, 284.4375, 284.4622, 284.4651, 
    284.4407, 284.4321, 284.321, 284.3083, 284.2036, 284.4573, 284.76, 
    278.1985, 281.5754, 286.355, 284.4695, 284.2446, 285.8481, 284.5208, 
    284.0386, 283.7251, 283.5264, 283.4595, 283.5212, 283.7937, 284.4019, 
    284.9829, 284.4617, 284.7075, 284.6848, 284.3792,
  282.2856, 281.9468, 281.6326, 281.575, 281.4634, 281.3926, 281.458, 
    281.4626, 281.5552, 281.1699, 281.1858, 281.7603, 281.5413, 281.4597, 
    280.7871, 280.7119, 280.9314, 280.6934, 280.7261, 280.7739, 282.521, 
    283.1333, 283.1133, 283.0706, 283.012, 282.6819, 282.5342, 282.5229, 
    282.5522, 282.6465, 282.8152, 282.939, 283.01, 283.0945, 283.2468, 
    283.3379, 283.4929, 284.043, 284.8599, 285.937, 286.5435, 285.3979, 
    285.5537, 285.5903, 285.9644, 279.7017, 286.2856, 286.9519, 286.843, 
    287.0083, 286.5137, 285.8088, 285.887, 285.603, 285.0356, 284.626, 
    284.3601, 284.0952, 283.9121, 283.7639, 283.6768, 283.5933, 283.3972, 
    283.2969, 283.1899, 283.0828, 283.0139, 282.917, 282.917, 282.8525, 
    282.9036, 282.946, 282.8921, 282.9285, 282.8743, 283.1362, 283.5342, 
    277.178, 282.2729, 285.3286, 282.2698, 281.3621, 281.8062, 281.885, 
    281.8479, 281.7383, 281.605, 281.4849, 281.5139, 281.4819, 281.804, 
    282.3257, 282.1604, 282.3794, 282.7297, 282.7644,
  280.1917, 280.1477, 279.9556, 279.9966, 279.875, 279.7637, 279.7554, 
    279.7124, 279.9998, 279.9233, 279.6924, 279.6809, 279.6687, 279.812, 
    279.4771, 279.2063, 279.3149, 278.7236, 279.2629, 279.0046, 280.4937, 
    281.1899, 281.1277, 281.0813, 281.0872, 280.9351, 280.6765, 280.5176, 
    280.4937, 280.5483, 280.7139, 280.9363, 281.1929, 281.3127, 281.6392, 
    282.0491, 282.0593, 282.4448, 282.8142, 283.1553, 283.3701, 283.2227, 
    283.3904, 283.5352, 284.106, 283.9807, 282.9712, 282.573, 282.3562, 
    282.6633, 282.5581, 282.3445, 282.7341, 283.4297, 283.2744, 282.8381, 
    282.6003, 282.3857, 282.2776, 282.187, 282.2168, 282.2734, 282.1475, 
    282.0513, 281.9395, 281.8545, 281.7373, 281.6118, 281.5693, 281.4502, 
    281.5444, 281.6211, 281.6272, 281.6985, 281.7244, 281.9675, 282.2861, 
    275.5303, 280.9338, 282.9224, 281.2041, 279.8354, 279.8052, 280.2192, 
    280.2036, 280.042, 280.0396, 279.9573, 280.0527, 280.0164, 280.0801, 
    280.1553, 280.2278, 280.2576, 280.1667, 280.4023,
  277.7578, 278.0688, 278.2686, 278.3259, 278.2395, 278.1968, 278.1763, 
    278.0962, 278.2605, 278.2634, 278.1809, 278.1533, 278.2661, 278.3108, 
    278.1467, 278.0676, 277.9497, 277.5669, 277.8071, 277.3879, 277.5293, 
    278.8694, 279.6692, 279.1838, 278.991, 278.8411, 278.7317, 278.6648, 
    278.6736, 278.7292, 278.8057, 278.9639, 279.2363, 279.3472, 279.5771, 
    280.311, 280.4368, 280.6025, 280.9744, 281.5498, 281.6179, 281.592, 
    281.8423, 281.895, 282.3362, 282.2324, 281.4856, 280.5186, 280.3188, 
    280.3921, 280.4468, 280.4089, 280.6821, 281.469, 281.5691, 281.355, 
    281.1416, 280.8184, 280.6511, 280.5708, 280.6707, 280.8728, 280.9104, 
    280.8455, 280.7561, 280.7549, 280.6545, 280.5225, 280.4282, 280.3022, 
    280.3464, 280.4163, 280.4338, 280.5381, 280.6531, 280.9321, 281.333, 
    276.135, 282.1904, 281.7471, 281.145, 279.8586, 278.9312, 278.8257, 
    278.6826, 278.3918, 278.489, 278.5625, 278.8401, 278.7756, 278.8384, 
    278.7212, 278.6628, 278.405, 277.5029, 277.7722,
  276.2527, 276.3787, 276.5828, 276.71, 276.7275, 276.7593, 276.7847, 
    276.7964, 276.7996, 276.8193, 276.9702, 276.9661, 277.0325, 277.0337, 
    276.9597, 276.9448, 276.8657, 276.5879, 276.3916, 275.9163, 275.4036, 
    274.627, 275.5752, 275.2961, 275.5503, 275.7092, 275.8872, 276.0869, 
    276.2747, 276.5288, 276.7402, 276.9519, 277.187, 277.3362, 277.5244, 
    278.0959, 278.4124, 278.4941, 278.3677, 278.9905, 279.3997, 279.4487, 
    280.0391, 280.2637, 280.9185, 281.4106, 280.7188, 279.0894, 278.8132, 
    278.8547, 278.8809, 279.0566, 279.5923, 279.8784, 279.7727, 279.6123, 
    279.4199, 279.0562, 279.0227, 278.9502, 279.1392, 279.3311, 279.5425, 
    279.5842, 279.4268, 279.5591, 279.5962, 279.5391, 279.4646, 279.3606, 
    279.335, 279.345, 279.3398, 279.394, 279.5129, 279.8174, 280.4133, 
    276.6123, 280.4717, 280.2322, 279.8928, 279.0552, 278.3528, 277.9478, 
    277.6633, 277.3726, 277.4192, 277.6353, 277.8479, 277.8096, 277.9177, 
    277.5969, 277.271, 276.9053, 276.2124, 276.2446,
  275.073, 274.9602, 274.8965, 275.1653, 275.311, 275.3586, 275.4097, 
    275.4963, 275.5554, 275.6113, 275.8081, 275.835, 275.8257, 275.8711, 
    275.8306, 275.7937, 275.7273, 275.5947, 275.3442, 274.4941, 273.8501, 
    273.0967, 272.8462, 272.5566, 272.6887, 272.9844, 273.261, 273.521, 
    273.8052, 274.1963, 274.5901, 274.9661, 275.2825, 275.5195, 275.739, 
    276.0625, 276.3855, 276.6353, 276.4961, 276.3511, 276.5737, 276.9678, 
    277.4668, 277.8391, 278.5366, 278.8003, 278.2354, 277.5769, 277.6443, 
    277.6694, 277.8438, 278.1233, 278.2483, 278.0823, 277.9045, 277.636, 
    277.0637, 276.7786, 277.4534, 277.4048, 277.4004, 277.4741, 277.7571, 
    277.991, 277.8643, 277.9778, 278.1257, 278.1533, 278.1726, 278.1401, 
    278.1746, 278.2092, 278.2317, 278.2456, 278.3215, 278.458, 279.0625, 
    279.5439, 276.0518, 279.1492, 278.5012, 277.9702, 277.5696, 277.4221, 
    277.2488, 276.8491, 276.573, 276.6821, 276.9629, 276.8948, 276.906, 
    276.5491, 276.2573, 276.0901, 275.6675, 275.3152,
  274.2039, 274.0005, 273.8501, 274.0164, 274.0713, 274.0322, 274.0608, 
    274.1882, 274.2737, 274.3384, 274.4597, 274.5481, 274.5974, 274.6165, 
    274.5732, 274.5005, 274.3845, 274.2795, 273.9841, 272.7642, 271.4646, 
    270.8938, 269.6931, 269.0249, 269.5647, 269.9529, 270.4067, 270.8469, 
    271.4001, 272.0254, 272.5608, 272.9978, 273.395, 273.7451, 274.0281, 
    274.3347, 274.6536, 274.8779, 274.9441, 274.8052, 274.9438, 275.3608, 
    275.8442, 276.4138, 276.8782, 276.772, 276.615, 276.6023, 276.6445, 
    276.6414, 276.6807, 276.6328, 276.5303, 276.137, 275.6592, 275.3279, 
    274.8928, 274.957, 276.0049, 276.0767, 275.9614, 276.0518, 276.2056, 
    276.3289, 276.364, 276.45, 276.5669, 276.6394, 276.6875, 276.7466, 
    276.7864, 276.874, 276.906, 276.958, 277.0183, 277.1343, 277.2725, 
    277.8289, 277.9788, 277.0957, 275.9797, 275.5437, 275.196, 275.5815, 
    275.6406, 275.5811, 275.4404, 275.4202, 275.7397, 275.6743, 275.6394, 
    275.1985, 274.9277, 274.8679, 274.8379, 274.5574,
  272.8662, 272.7241, 272.6077, 272.6445, 272.6736, 272.697, 272.7346, 
    272.8169, 272.8779, 272.9104, 272.9604, 273.0757, 273.1555, 273.1326, 
    273.0134, 272.8193, 272.6318, 272.4822, 272.2783, 271.0537, 268.9036, 
    268.2307, 266.8606, 265.7961, 266.512, 267.1331, 267.6543, 268.2546, 
    268.9736, 269.6777, 270.3967, 271.0552, 271.6143, 272.0803, 272.4385, 
    272.7258, 272.7041, 272.9016, 272.9951, 273.0515, 273.3027, 273.5178, 
    273.7908, 274.238, 274.4368, 274.4126, 274.6733, 274.9314, 274.9556, 
    274.8237, 274.5439, 274.1875, 274.1121, 273.7893, 273.2488, 273.1538, 
    273.3743, 273.8171, 274.3765, 274.3164, 274.3394, 274.575, 274.6904, 
    274.8474, 274.9822, 275.0874, 275.1865, 275.2712, 275.3352, 275.4104, 
    275.4636, 275.5078, 275.5535, 275.5989, 275.6653, 275.7292, 275.7012, 
    275.7327, 275.2385, 274.3157, 273.7883, 273.3577, 273.0186, 273.1343, 
    273.4783, 273.6113, 273.7351, 273.8716, 273.98, 273.9041, 273.728, 
    273.259, 273.0659, 273.1519, 273.2795, 273.0974,
  271.0723, 270.8071, 270.6455, 270.7976, 270.8359, 270.9238, 271.0806, 
    271.2451, 271.2175, 271.1106, 271.1384, 271.3037, 271.2075, 270.7026, 
    269.9622, 268.9949, 268.4043, 268.1116, 267.8745, 266.9929, 265.4592, 
    264.8125, 263.7673, 262.8374, 263.4097, 263.9844, 264.2334, 264.3772, 
    264.843, 265.6987, 266.4224, 267.0283, 267.9253, 268.6743, 269.1758, 
    269.2346, 268.8535, 269.0283, 268.8457, 269.0586, 269.8115, 270.2065, 
    270.4346, 270.8003, 271.1909, 271.3633, 271.6694, 272.0015, 271.9602, 
    271.7329, 271.541, 271.1558, 271.0742, 270.9382, 270.7417, 271.2874, 
    271.905, 272.2668, 272.3494, 272.2515, 272.4314, 272.6943, 272.9065, 
    273.1743, 273.3196, 273.4282, 273.5632, 273.6846, 273.7874, 273.9319, 
    274.0442, 274.1174, 274.2456, 274.332, 274.376, 274.3594, 274.2202, 
    273.948, 273.4966, 272.3052, 270.675, 270.1924, 269.7859, 270.3296, 
    270.9448, 271.0476, 271.303, 271.5464, 271.6348, 271.687, 271.4121, 
    270.9326, 271.2278, 271.6387, 271.6831, 271.3403,
  268.4519, 268.2466, 268.0649, 267.9678, 267.7773, 268.0181, 268.3745, 
    268.5776, 267.8145, 267.45, 267.6636, 267.4375, 265.5415, 262.2861, 
    260.6201, 259.5098, 258.9653, 259.4575, 260.0261, 260.4172, 260.1331, 
    259.7913, 259.7092, 258.2222, 258.8557, 259.2747, 259.3, 259.4497, 
    259.6965, 259.8271, 260.0046, 260.415, 261.061, 261.4446, 261.6323, 
    261.3848, 260.7644, 260.2708, 259.8279, 260.9458, 262.6519, 263.2913, 
    263.5657, 264.4524, 265.5312, 266.1409, 266.905, 267.5168, 267.5781, 
    267.4326, 267.7817, 267.7937, 267.793, 268.0527, 268.8789, 269.7659, 
    270.2937, 270.1409, 269.7305, 269.8721, 270.2708, 270.4473, 270.5984, 
    270.8572, 271.0808, 271.3347, 271.595, 271.8403, 272.1211, 272.4177, 
    272.6653, 272.8853, 273.0806, 273.157, 273.2109, 273.2058, 273.0588, 
    272.6748, 271.9521, 264.8176, 267.4438, 267.3127, 267.5347, 267.9519, 
    268.217, 268.1021, 268.2505, 268.4521, 268.5393, 268.3318, 267.988, 
    268.1155, 268.7031, 268.7861, 268.6035, 268.4983,
  264.8467, 264.5129, 264.2554, 263.6985, 262.9517, 262.8083, 262.8621, 
    263.2488, 260.9753, 261.6047, 262.1321, 262.196, 262.8381, 251.0445, 
    251.4453, 249.9639, 255.2595, 255.5579, 255.1525, 255.5599, 256.0522, 
    256.9841, 259.4343, 251.9276, 250.1555, 249.1581, 248.5105, 247.647, 
    247.9915, 249.7699, 250.8578, 252.3495, 252.952, 252.7107, 251.3766, 
    248.8177, 247.3784, 248.3781, 250.5004, 256.4438, 257.5347, 256.5759, 
    256.0098, 257.2979, 258.6968, 259.9407, 261.6897, 262.7915, 263.2578, 
    263.5461, 263.9583, 264.0632, 264.4126, 265.1877, 266.1768, 266.9504, 
    267.282, 267.0515, 266.8562, 267.0703, 267.3188, 267.4211, 267.5889, 
    268.0002, 268.4963, 269.0044, 269.4851, 269.96, 270.4629, 270.9387, 
    271.2437, 271.427, 271.5842, 271.7139, 271.9377, 272.0576, 271.6292, 
    270.2825, 261.3369, 261.0127, 264.5205, 264.5842, 265.2078, 265.6311, 
    265.6899, 265.4675, 265.3887, 265.3992, 265.3057, 265.1152, 265.0317, 
    265.0215, 264.9895, 264.8835, 265.0144, 265.0547,
  259.6206, 259.927, 260.1318, 260.1086, 259.8049, 259.7563, 260.2461, 
    263.1748, 251.1971, 255.1997, 253.1543, 249.9514, 245.5794, 243.1769, 
    238.8615, 236.2359, 240.6458, 243.1568, 244.2042, 244.3191, 249.4648, 
    249.0741, 244.8095, 239.518, 236.901, 236.1926, 235.89, 236.1945, 
    237.1453, 238.4371, 239.4215, 240.276, 240.6164, 239.5273, 237.767, 
    236.0851, 236.8085, 238.2018, 241.3891, 242.6696, 245.0865, 246.7194, 
    247.3197, 252.7767, 252.1139, 252.6588, 255.3168, 257.1497, 258.3013, 
    258.9988, 259.5835, 260.177, 261.001, 261.9355, 262.7017, 263.177, 
    263.4397, 263.5535, 263.772, 264.0762, 264.1133, 264.343, 264.708, 
    265.2734, 265.9258, 266.512, 267.051, 267.5933, 268.2671, 268.6489, 
    268.8613, 268.9307, 269.2163, 269.5984, 270.2522, 270.7944, 270.5884, 
    258.9075, 258.4583, 257.1472, 260.8523, 261.5598, 262.4634, 263.0068, 
    262.9602, 262.6633, 262.4395, 262.3113, 262.0996, 261.7598, 261.1135, 
    260.54, 260.0535, 258.6458, 258.925, 259.3169,
  246.4325, 242.8583, 239.4129, 237.2406, 238.0668, 240.7682, 241.1096, 
    239.9867, 239.0478, 237.9484, 236.8074, 233.5639, 229.5863, 226.7626, 
    226.5911, 229.7815, 232.767, 234.4168, 234.8202, 240.279, 242.6341, 
    240.0539, 232.9902, 227.1163, 225.9549, 226.1562, 226.7329, 226.9344, 
    227.3306, 227.0977, 227.4941, 227.9526, 227.528, 227.0658, 227.5316, 
    228.0891, 228.9396, 229.1341, 229.4875, 231.8382, 233.6876, 236.0614, 
    239.1745, 242.0273, 244.0562, 249.6484, 251.6967, 252.9536, 254.1224, 
    255.2236, 256.1047, 256.7446, 257.3506, 258.0276, 258.8086, 259.5391, 
    260.0176, 260.2402, 260.5129, 261.2229, 260.9744, 261.3801, 261.6714, 
    261.9646, 262.5435, 262.8774, 263.3206, 263.686, 264.1035, 264.5503, 
    264.6736, 264.8315, 264.8965, 264.9709, 265.6106, 266.4209, 266.1672, 
    253.6879, 255.0036, 255.0842, 257.1245, 258.4033, 259.3933, 259.9172, 
    259.9412, 259.7114, 259.4285, 259.0798, 258.7539, 258.0938, 256.9001, 
    257.3862, 260.1101, 251.1825, 250.9267, 248.5602,
  230.7305, 227.918, 226.2072, 225.0434, 224.8497, 225.0387, 224.3789, 
    223.7048, 223.1069, 223.1917, 223.6915, 223.8388, 223.6895, 224.0165, 
    226.5025, 229.0698, 230.7238, 232.593, 234.9583, 235.6017, 237.3501, 
    231.7324, 228.1594, 224.0296, 221.3421, 219.6523, 219.4085, 219.9941, 
    220.54, 221.297, 221.1232, 220.7121, 220.6215, 220.9133, 222.082, 
    223.8176, 225.2844, 226.2599, 227.2186, 229.0053, 231.3961, 235.0159, 
    238.7477, 243.8361, 243.6839, 250.1495, 250.7298, 250.6943, 250.8872, 
    251.8976, 252.8559, 253.5413, 254.1073, 254.6279, 255.3008, 256.1089, 
    256.574, 257.1104, 257.948, 259.7327, 252.3301, 253.0725, 253.0233, 
    253.1686, 253.3204, 253.1295, 253.4729, 254.4624, 255.1569, 254.5546, 
    253.7272, 251.445, 248.8215, 247.9208, 248.5087, 249.7026, 250.3249, 
    250.0736, 250.7613, 248.6323, 254.0717, 255.2618, 256.2681, 256.6633, 
    256.7271, 256.6162, 256.6123, 256.2456, 255.7605, 257.6431, 252.3156, 
    250.638, 245.3762, 241.8246, 237.2159, 233.4782,
  225.6796, 223.5928, 220.9743, 218.5699, 218.0535, 217.8102, 217.3427, 
    217.1117, 217.0284, 217.5958, 218.1361, 219.3529, 220.9346, 222.6476, 
    224.5979, 226.7348, 229.12, 230.0133, 229.9193, 229.1811, 227.1561, 
    224.8559, 221.979, 218.9331, 217.5794, 216.7194, 216.9105, 217.8073, 
    218.4456, 218.5788, 218.7314, 218.9741, 219.4622, 220.5883, 222.7958, 
    224.3596, 225.3436, 226.0299, 227.2311, 228.7979, 231.463, 234.8927, 
    239.4018, 246.1251, 247.5423, 247.2586, 245.3077, 243.6678, 242.8458, 
    242.9633, 243.5598, 244.3382, 245.129, 246.3798, 247.5621, 248.6275, 
    249.8021, 251.1016, 251.9874, 250.3612, 248.4523, 247.0539, 246.3289, 
    246.2279, 246.5077, 246.8501, 247.8902, 248.6264, 248.8566, 248.4734, 
    246.901, 245.318, 245.6555, 246.594, 246.381, 247.1219, 246.5855, 
    245.966, 245.4005, 245.5775, 251.1088, 252.4325, 253.2366, 253.7066, 
    253.925, 253.8579, 254.2031, 255.56, 251.1409, 251.1724, 247.3978, 
    242.424, 237.5435, 232.4469, 228.843, 226.9449,
  226.6168, 225.2701, 223.138, 221.8025, 220.7126, 219.3581, 217.8335, 
    216.849, 216.722, 216.2086, 216.1752, 216.4125, 216.7441, 217.4115, 
    217.6078, 217.9499, 218.3301, 218.8302, 218.9921, 218.0651, 217.4426, 
    216.3578, 215.2833, 214.7467, 213.9017, 214.4252, 215.3387, 217.0552, 
    218.8134, 219.3868, 219.6654, 220.0099, 220.6927, 223.431, 225.2436, 
    226.453, 227.1012, 228.7667, 230.1557, 232.6715, 236.5375, 240.0988, 
    244.2139, 246.0795, 245.9797, 246.2137, 245.8874, 244.8272, 244.1555, 
    243.7975, 243.5401, 243.4215, 244.1139, 244.7134, 244.7449, 245.0207, 
    245.8251, 246.7184, 246.6256, 247.1969, 247.5383, 247.3371, 247.0226, 
    246.2906, 245.2577, 245.0807, 244.4657, 243.3062, 241.9838, 240.8962, 
    240.4325, 241.0215, 242.854, 245.6913, 247.8432, 248.1696, 246.9642, 
    245.1772, 243.5668, 243.6717, 244.0603, 243.7393, 243.9885, 244.5048, 
    245.7398, 247.8867, 249.9264, 251.6151, 250.8532, 250.3949, 246.2521, 
    240.4255, 235.9379, 230.6415, 227.7358, 227.2952,
  229.0755, 227.8814, 226.5146, 224.3546, 222.5109, 221.1292, 220.1087, 
    219.022, 217.8708, 216.7421, 215.797, 215.0595, 214.6926, 214.3719, 
    214.187, 213.9927, 213.8326, 213.3068, 212.978, 212.8002, 212.6668, 
    213.501, 214.3216, 214.6483, 215.7227, 216.2577, 217.7828, 219.1863, 
    220.6289, 221.4905, 221.666, 222.5237, 223.6224, 225.3825, 227.1195, 
    227.5838, 228.923, 231.056, 232.526, 234.8948, 237.5288, 239.501, 
    242.4471, 246.9622, 249.8029, 249.9476, 249.6952, 249.5883, 249.0078, 
    248.1887, 247.2914, 246.1443, 245.1009, 244.5589, 244.1355, 243.6423, 
    242.7609, 242.7379, 243.287, 244.3758, 245.7414, 247.518, 248.9974, 
    249.832, 249.1737, 247.2005, 244.5453, 241.2444, 239.848, 238.5909, 
    237.5422, 237.6928, 239.0169, 241.5381, 243.1881, 245.0264, 245.6178, 
    246.2101, 246.4749, 246.409, 247.2798, 247.5509, 247.3268, 247.8324, 
    249.4605, 251.1333, 249.5565, 247.5465, 245.8531, 244.1181, 241.0023, 
    237.2079, 234.387, 230.8973, 229.5943, 229.5924,
  226.6716, 226.6732, 226.335, 224.0323, 224.21, 224.1893, 224.1672, 
    223.9611, 223.3146, 222.6371, 221.9688, 221.341, 220.4471, 219.7045, 
    219.2087, 218.3615, 217.5237, 216.7405, 216.4297, 216.5484, 216.8441, 
    217.9944, 218.629, 219.1191, 219.3647, 219.6424, 220.0074, 220.643, 
    221.2406, 221.937, 222.6499, 223.3991, 223.9543, 224.8936, 226.0936, 
    226.4144, 226.425, 228.4122, 230.2421, 231.706, 232.424, 232.4469, 
    235.1483, 237.1629, 238.4264, 239.2923, 239.9958, 241.8272, 244.8233, 
    247.0033, 248.1263, 249.244, 249.6411, 250.0036, 250.4637, 250.1075, 
    249.6046, 249.4229, 249.0766, 248.3975, 247.3236, 246.1746, 245.2798, 
    244.0961, 242.2988, 240.5462, 238.2715, 236.0984, 235.0487, 233.8811, 
    234.1625, 234.6109, 235.6174, 237.5819, 240.1448, 241.9165, 243.4997, 
    244.1495, 244.7902, 245.0522, 244.9874, 244.6605, 243.7809, 243.1405, 
    242.5363, 241.2353, 239.8284, 238.4799, 237.1381, 235.4915, 233.634, 
    232.3956, 230.4501, 228.7625, 227.8102, 227.0118,
  225.8387, 225.7345, 226.1768, 225.8551, 225.6023, 225.5207, 225.4151, 
    225.3792, 225.5609, 225.4782, 225.0389, 224.1358, 223.224, 222.6621, 
    222.6392, 222.7478, 222.7566, 222.4932, 222.0631, 221.9107, 221.5475, 
    221.5066, 221.7038, 221.5448, 221.578, 221.8051, 221.6732, 222.1395, 
    222.2643, 222.4262, 222.1978, 222.2377, 222.4025, 223.1387, 223.8961, 
    224.1083, 224.1905, 224.2366, 224.3181, 224.4891, 224.95, 225.5178, 
    226.147, 226.7914, 228.1139, 229.5134, 229.8519, 229.6453, 229.0488, 
    228.7188, 229.2747, 230.0335, 230.6104, 231.4393, 232.3181, 233.1026, 
    233.8543, 234.3763, 234.7553, 235.2828, 235.6737, 236.1453, 236.2228, 
    235.9362, 235.6169, 235.419, 235.3151, 235.1004, 235.2234, 235.6767, 
    235.8424, 236.0651, 237.0759, 238.0849, 238.1372, 237.4034, 236.3419, 
    234.9406, 233.7858, 233.0042, 232.5056, 232.2137, 232.3831, 232.1715, 
    232.4682, 231.1848, 230.0684, 229.5751, 228.4039, 228.642, 228.6684, 
    228.3083, 227.1579, 226.7548, 226.5596, 226.0381,
  228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 
    228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 
    228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 
    228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 
    228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 
    228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 
    228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 
    228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 
    228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 
    228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 
    228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 
    228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 
    228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 228.4698, 
    228.4698, 228.4698, 228.4698, 228.4698, 228.4698 ;
}
